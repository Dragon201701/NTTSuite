
--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/ccs_libs/interfaces/amba/amba_comps.vhd 
--//////////////////////////////////////////////////////////////////////////////
-- Catapult Synthesis - Custom Interfaces
--
-- Copyright (c) 2016 Mentor Graphics Corp.
--       All Rights Reserved
-- 
-- This document contains information that is proprietary to Mentor Graphics
-- Corp. The original recipient of this document may duplicate this  
-- document in whole or in part for internal business purposes only, provided  
-- that this entire notice appears in all copies. In duplicating any part of  
-- this document, the recipient agrees to make every reasonable effort to  
-- prevent the unauthorized use and distribution of the proprietary information.
-- 
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in prepartion for creating
-- their own custom interfaces. This design does not present a complete
-- implementation of the named protocol or standard.
--
-- NO WARRANTY.
-- MENTOR GRAPHICS CORP. EXPRESSLY DISCLAIMS ALL WARRANTY
-- FOR THE SOFTWARE. TO THE MAXIMUM EXTENT PERMITTED BY APPLICABLE
-- LAW, THE SOFTWARE AND ANY RELATED DOCUMENTATION IS PROVIDED "AS IS"
-- AND WITH ALL FAULTS AND WITHOUT WARRANTIES OR CONDITIONS OF ANY
-- KIND, EITHER EXPRESS OR IMPLIED, INCLUDING, WITHOUT LIMITATION, THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR
-- PURPOSE, OR NONINFRINGEMENT. THE ENTIRE RISK ARISING OUT OF USE OR
-- DISTRIBUTION OF THE SOFTWARE REMAINS WITH YOU.
-- 
--//////////////////////////////////////////////////////////////////////////////

-- --------------------------------------------------------------------------
-- LIBRARY: amba
--
-- CONTENTS:
--    axi4stream_w_wire, axi4stream_r_wire, axi4svideo_w_wire, axi4svideo_r_wire
--      Catapult AXI-4 Stream bus definitions
--    ccs_axi4stream_in
--      AXI4-Streaming input interface
--    ccs_axi4stream_out
--      AXI4-Streaming output interface
--    ccs_axi4stream_pipe
--      AXI4-Streaming FIFO interconnect component
--    ccs_axi4svideo_in
--      AXI4-Streaming video input interface
--    ccs_axi4svideo_out
--      AXI4-Streaming video output interface
--    ccs_axi4svideo_pipe
--      AXI4-Streaming video FIFO interconnect component
--
--    axi4_busdef
--      Catapult AXI-4 bus definition
--
--    ccs_axi4_slave_mem
--      Catapult AXI-4 slave memory
---
--    ccs_axi4_master
--      Catapult AXI4 master interface for read/write data
--
--    apb_busdef
--      Catapult APB bus definition
--    apb_slave_mem
--      APB Slave Memory interface
--
-- CHANGE LOG:
--
--  10/01/16 - dgb - Initial implementation
--
-- --------------------------------------------------------------------------

-- --------------------------------------------------------------------------
-- PACKAGE:     amba_comps
--
-- DESCRIPTION:
--   Contains component declarations for all design units in this file.
--
-- CHANGE LOG:
--
--  10/01/16 - dgb - Initial implementation
--
-- --------------------------------------------------------------------------

LIBRARY ieee;

   USE ieee.std_logic_1164.all;
   USE ieee.std_logic_arith.all;
   USE ieee.std_logic_unsigned.all;

PACKAGE amba_comps IS

  -- ==============================================================
  -- AXI-4 Stream Components
  -- ------------------------------ TSTRB/TKEEP controls --------------------
  --    TKEEP   TSTRB   Data Type         Description
  --    high    high    Data byte         Valid data byte (supported in these models)
  --    high    low     Position byte     Byte is position not data/null (not supported)
  --    low     low     Null byte         Byte is null (not supported)
  --    low     high    Reserved          Do not use (not supported)

  COMPONENT axi4stream_w_wire -- slave interface pin direction
    GENERIC(
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 16;           -- AXI4 Bus width
      AXI4_USER_WIDTH  : INTEGER RANGE 1 TO 8 := 1                -- AXI4 User data width
    );
    PORT(
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : IN   std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : OUT  std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : IN   std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TLAST     : IN   std_logic;                                        -- M->S      Indicates boundary of a packet
      TUSER     : IN   std_logic_vector(AXI4_USER_WIDTH-1 downto 0)      -- M->S      Optional user-defined sideband data
    );
  END COMPONENT;

  COMPONENT axi4stream_r_wire -- master interface pin direction
    GENERIC(
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 16;           -- AXI4 Bus width
      AXI4_USER_WIDTH  : INTEGER RANGE 1 TO 8 := 1                -- AXI4 User data width
    );
    PORT(
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : OUT  std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : IN   std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : OUT  std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TLAST     : OUT  std_logic;                                        -- M->S      Indicates boundary of a packet
      TUSER     : OUT  std_logic_vector(AXI4_USER_WIDTH-1 downto 0)      -- M->S      Optional user-defined sideband data
    );
  END COMPONENT;

  COMPONENT axi4svideo_w_wire -- slave interface pin direction
    GENERIC(
      width            : INTEGER RANGE 3 TO 1024 := 33;           -- Catapult read/write operator width
      AXI4_DATA_WIDTH  : INTEGER                 := 16            -- AXI4 Bus width
    );
    PORT(
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : IN   std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : OUT  std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : IN   std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TUSER     : IN   std_logic;                                        -- M->S      Start of Frame
      TLAST     : IN   std_logic                                         -- M->S      End of Line
    );
  END COMPONENT;

  COMPONENT axi4svideo_r_wire -- master interface pin direction
    GENERIC(
      width            : INTEGER RANGE 3 TO 1024 := 33;           -- Catapult read/write operator width
      AXI4_DATA_WIDTH  : INTEGER                 := 16            -- AXI4 Bus width
    );
    PORT(
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : OUT  std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : IN   std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : OUT  std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TUSER     : OUT  std_logic;                                        -- M->S      Start of Frame
      TLAST     : OUT  std_logic                                         -- M->S      End of Line
    );
  END COMPONENT;

  COMPONENT ccs_axi4stream_in
    GENERIC(
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 32;           -- AXI4 Bus width
      AXI4_USER_WIDTH  : INTEGER RANGE 1 TO 8 := 1                -- AXI4 User data width
    );
    PORT(
      -- AXI-4 Master Clock/Reset
      ACLK      : IN   std_logic;                                        -- clk src   Rising edge clock
      ARESETn   : IN   std_logic;                                        -- rst src   Active LOW synchronous reset
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : IN   std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : OUT  std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : IN   std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TLAST     : IN   std_logic;                                        -- M->S      Indicates boundary of a packet
      TUSER     : IN   std_logic_vector(AXI4_USER_WIDTH-1 downto 0);     -- M->S      Optional user-defined sideband data
      -- Catapult interface (equiv to mgc_in_wire_wait)
      d         : OUT  std_logic_vector(width-1 downto 0);               -- d  - msb TLAST TUSER(...) TDATA(...) lsb
      vd        : OUT  std_logic;                                        -- vd - TVALID
      ld        : IN   std_logic                                         -- ld - TREADY
    );
  END COMPONENT;

  COMPONENT ccs_axi4stream_out
    GENERIC(
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 32;           -- AXI4 Bus width
      AXI4_USER_WIDTH  : INTEGER RANGE 1 TO 8 := 1                -- AXI4 User data width
    );
    PORT(
      -- AXI-4 Master Clock/Reset
      ACLK      : IN   std_logic;                                        -- clk src   Rising edge clock
      ARESETn   : IN   std_logic;                                        -- rst src   Active LOW synchronous reset
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : OUT  std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : IN   std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : OUT  std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TLAST     : OUT  std_logic;                                        -- M->S      Indicates boundary of a packet
      TUSER     : OUT  std_logic_vector(AXI4_USER_WIDTH-1 downto 0);     -- M->S      Optional user-defined sideband data
      -- Catapult interface (equiv to mgc_out_stdreg_wait)
      d         : IN   std_logic_vector(width-1 downto 0);               -- d  - msb TLAST TUSER(...) TDATA(...) lsb
      vd        : OUT  std_logic;                                        -- vd - TREADY
      ld        : IN   std_logic                                         -- ld - TVALID
    );
  END COMPONENT;

  -- This implementation currently does not work - the 'width' parameter is not configured properly
  COMPONENT ccs_axi4stream_pipe
    GENERIC(
      rscid            : INTEGER := 1;                            -- Resource ID from Catapult
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      fifo_sz          : INTEGER RANGE 0 TO 128 := 0;            -- Fifo size
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 32;           -- AXI4 Bus width
      AXI4_USER_WIDTH  : INTEGER RANGE 1 TO 8 := 1                -- AXI4 User data width
    );
    PORT(
      -- AXI-4 Master Clock/Reset
      ACLK      : IN   std_logic;                                          -- clk src   Rising edge clock
      ARESETn   : IN   std_logic;                                          -- rst src   Active LOW asynchronous reset
      -- AXI-4 Stream interface input                                      -- Src->Dst  Description
      sTVALID   : IN   std_logic;                                          -- M->S      Indicates master is driving a valid transfer
      sTREADY   : OUT  std_logic;                                          -- S->M      Indicates slave can accept a transfer
      sTDATA    : IN   std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);       -- M->S      Primary payload (width-1 must be multiple of 8)
      sTSTRB    : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 indicates data byte, 0 indicates position byte
      sTKEEP    : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 valid byte, 0 indicates null byte
      sTLAST    : IN   std_logic;                                          -- M->S      Indicates boundary of a packet
      sTUSER    : IN   std_logic_vector(AXI4_USER_WIDTH-1 downto 0);       -- M->S      Optional user-defined sideband data
      -- AXI-4 Stream interface output                                     -- Src->Dst  Description
      mTVALID   : OUT  std_logic;                                          -- M->S      Indicates master is driving a valid transfer
      mTREADY   : IN   std_logic;                                          -- S->M      Indicates slave can accept a transfer
      mTDATA    : OUT  std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);       -- M->S      Primary payload (width-1 must be multiple of 8)
      mTSTRB    : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 indicates data byte, 0 indicates position byte
      mTKEEP    : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 valid byte, 0 indicates null byte
      mTLAST    : OUT  std_logic;                                          -- M->S      Indicates boundary of a packet
      mTUSER    : OUT  std_logic_vector(AXI4_USER_WIDTH-1 downto 0)        -- M->S      Optional user-defined sideband data
    );
  END COMPONENT;

  COMPONENT ccs_axi4svideo_in
    GENERIC(
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 32            -- AXI4 Bus width
    );
    PORT(
      -- AXI-4 Master Clock/Reset
      ACLK      : IN   std_logic;                                        -- clk src   Rising edge clock
      ARESETn   : IN   std_logic;                                        -- rst src   Active LOW asynchronous reset
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : IN   std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : OUT  std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : IN   std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TLAST     : IN   std_logic;                                        -- M->S      End-of-line
      TUSER     : IN   std_logic;                                        -- M->S      Start-of-frame
      -- Catapult interface (equiv to mgc_in_wire_wait)
      d         : OUT  std_logic_vector(width-1 downto 0);               -- d  - msb TLAST TUSER TDATA(...) lsb
      vd        : OUT  std_logic;                                        -- vd - TVALID
      ld        : IN   std_logic                                         -- ld - TREADY
    );
  END COMPONENT;

  COMPONENT ccs_axi4svideo_out
    GENERIC(
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 32            -- AXI4 Bus width
    );
    PORT(
      -- AXI-4 Master Clock/Reset
      ACLK      : IN   std_logic;                                        -- clk src   Rising edge clock
      ARESETn   : IN   std_logic;                                        -- rst src   Active LOW asynchronous reset
      -- AXI-4 Stream interface                                          -- Src->Dst  Description
      TVALID    : OUT  std_logic;                                        -- M->S      Indicates master is driving a valid transfer
      TREADY    : IN   std_logic;                                        -- S->M      Indicates slave can accept a transfer
      TDATA     : OUT  std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);     -- M->S      Primary payload (width-1 must be multiple of 8)
      TSTRB     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 indicates data byte, 0 indicates position byte
      TKEEP     : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0); -- M->S      1 valid byte, 0 indicates null byte
      TLAST     : OUT  std_logic;                                        -- M->S      End-of-line
      TUSER     : OUT  std_logic;                                        -- M->S      Start-of-frame
      -- Catapult interface (equiv to mgc_out_stdreg_wait)
      d         : IN   std_logic_vector(width-1 downto 0);               -- d  - msb TLAST TUSER TDATA(...) lsb
      vd        : OUT  std_logic;                                        -- vd - TREADY
      ld        : IN   std_logic                                         -- ld - TVALID
    );
  END COMPONENT;

  COMPONENT ccs_axi4svideo_pipe
    GENERIC(
      rscid            : INTEGER := 1;                                 -- Resource ID from Catapult
      width            : INTEGER RANGE 3 TO 1026 := 33;           -- Catapult read/write operator width (includes data,last and user bits)
      fifo_sz          : INTEGER RANGE 0 TO 128 := 0;            -- Fifo size
      AXI4_DATA_WIDTH  : INTEGER RANGE 8 TO 1024 := 32            -- AXI4 Bus width
    );
    PORT(
      -- AXI-4 Master Clock/Reset
      ACLK      : IN   std_logic;                                          -- clk src   Rising edge clock
      ARESETn   : IN   std_logic;                                          -- rst src   Active LOW asynchronous reset
      -- AXI-4 Stream interface input                                      -- Src->Dst  Description
      sTVALID   : IN   std_logic;                                          -- M->S      Indicates master is driving a valid transfer
      sTREADY   : OUT  std_logic;                                          -- S->M      Indicates slave can accept a transfer
      sTDATA    : IN   std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);       -- M->S      Primary payload (width-1 must be multiple of 8)
      sTSTRB    : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 indicates data byte, 0 indicates position byte
      sTKEEP    : IN   std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 valid byte, 0 indicates null byte
      sTLAST    : IN   std_logic;                                          -- M->S      End-of-line
      sTUSER    : IN   std_logic;                                          -- M->S      Start-of-frame
      -- AXI-4 Stream interface output                                     -- Src->Dst  Description
      mTVALID   : OUT  std_logic;                                          -- M->S      Indicates master is driving a valid transfer
      mTREADY   : IN   std_logic;                                          -- S->M      Indicates slave can accept a transfer
      mTDATA    : OUT  std_logic_vector(AXI4_DATA_WIDTH-1 downto 0);       -- M->S      Primary payload (width-1 must be multiple of 8)
      mTSTRB    : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 indicates data byte, 0 indicates position byte
      mTKEEP    : OUT  std_logic_vector((AXI4_DATA_WIDTH/8)-1 downto 0);   -- M->S      1 valid byte, 0 indicates null byte
      mTLAST    : OUT  std_logic;                                          -- M->S      End-of-line
      mTUSER    : OUT  std_logic                                           -- M->S      Start-of-frame
    );
  END COMPONENT;

  -- ==============================================================
  -- AXI-4 Bus Components

  -- Used to define the AXI-4 bus definition (direction of signals is from the slave's perspective)
    -- Pin directions are based on the usage of this busdef as a "master" driving an input slave.
    -- To use the bus in the reverse direction set the interface to "slave".
  COMPONENT axi4_busdef -- 
    GENERIC(   
      host_tidw      : INTEGER RANGE 1 TO 11 := 4;            -- Width of transaction ID fields
      host_userw     : INTEGER RANGE 1 TO 16 := 4;            -- Width of user-defined signals
      ADDR_WIDTH     : INTEGER RANGE 1 TO 64 := 32;           -- Host address width
      DATA_WIDTH     : INTEGER RANGE 8 TO 64 := 8             -- Host data width
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                 -- Rising edge clock
      ARESETn    : IN   std_logic;                                 -- Active LOW synchronous reset

      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(host_tidw-1 downto 0);    -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);      -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);              -- Write burst length    - must always be 0 in AXI4-Lite
      AWSIZE     : OUT  std_logic_vector(1 downto 0);              -- Write burst size      - must equal host_dw_bytes-2
      AWBURST    : OUT  std_logic_vector(1 downto 0);              -- Write burst mode      - must always be 0 (fixed mode) in AXI4-Lite
      AWLOCK     : OUT  std_logic;                                 -- Lock type             - must always be 0 (Normal access) in AXI4-Lite
      AWCACHE    : OUT  std_logic_vector(3 downto 0);              -- Memory type           - must always be 0 (Non-modifiable, Non-bufferable) in AXI4-Lite
      AWPROT     : OUT  std_logic_vector(2 downto 0);              -- Protection Type       - ignored in this model
      AWQOS      : OUT  std_logic_vector(3 downto 0);              -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);              -- Region identifier
      AWUSER     : OUT  std_logic_vector(host_userw-1 downto 0);   -- User signal
      AWVALID    : OUT  std_logic;                                 -- Write address valid
      AWREADY    : IN   std_logic;                                 -- Write address ready (slave is ready to accept AWADDR)
      
      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0); -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise) - ignored in AXI-4 Lite
      WLAST      : OUT  std_logic;                                        -- Write last
      WUSER      : OUT  std_logic_vector(host_userw-1 downto 0);          -- User signal
      WVALID     : OUT  std_logic;                                        -- Write data is valid
      WREADY     : IN   std_logic;                                        -- Write ready (slave is ready to accept WDATA)
      
      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(host_tidw-1 downto 0);    -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);              -- Write response (of slave) - only OKAY, SLVERR, DECERR supported in AXI-4 Lite
      BUSER      : IN   std_logic_vector(host_userw-1 downto 0);   -- User signal
      BVALID     : IN   std_logic;                                 -- Write response valid (slave accepted WDATA)
      BREADY     : OUT  std_logic;                                 -- Response ready (master can accept slave's write response)
      
      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(host_tidw-1 downto 0);    -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);      -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);              -- Read burst length     - must always be 0 in AXI4-Lite
      ARSIZE     : OUT  std_logic_vector(1 downto 0);              -- Read burst size       - must equal host_dw_bytes-2
      ARBURST    : OUT  std_logic_vector(1 downto 0);              -- Read burst mode       - must always be 0 (fixed mode) in AXI4-Lite
      ARLOCK     : OUT  std_logic;                                 -- Lock type             - must always be 0 (Normal access) in AXI4-Lite
      ARCACHE    : OUT  std_logic_vector(3 downto 0);              -- Memory type           - must always be 0 (Non-modifiable, Non-bufferable) in AXI4-Lite
      ARPROT     : OUT  std_logic_vector(2 downto 0);              -- Protection Type       - ignored in this model
      ARQOS      : OUT  std_logic_vector(3 downto 0);              -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);              -- Region identifier
      ARUSER     : OUT  std_logic_vector(host_userw-1 downto 0);   -- User signal
      ARVALID    : OUT  std_logic;                                 -- Read address valid
      ARREADY    : IN   std_logic;                                 -- Read address ready (slave is ready to accept ARADDR)
      
      -- ============== AXI4 Read Data Channel Signals
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0); -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                      -- Read response (of slave) - only OKAY, SLVERR, DECERR supported in AXI-4 Lite
      RVALID     : IN   std_logic;                                         -- Read valid (slave providing RDATA)
      RREADY     : OUT  std_logic;                                         -- Read ready (master ready to receive RDATA)
      RID        : OUT  std_logic_vector(host_tidw-1 downto 0);            -- Read ID tag
      RLAST      : IN   std_logic;                                         -- Read last
      RUSER      : IN   std_logic_vector(host_userw-1 downto 0)            -- User signal
    );
  END COMPONENT;

  -- AXI4 Lite GPIO with CDC
  COMPONENT ccs_axi4_lite_slave_cdc
    GENERIC(
      rscid          : INTEGER               := 1;            -- Required resource ID parameter
      op_width       : INTEGER RANGE 1 TO 64 := 1;            -- Operator width (dummy parameter)
      cwidth         : INTEGER RANGE 1 TO 256 := 32;          -- Internal register width
      nopreload      : INTEGER RANGE 0 TO 1 := 0;             -- 1=disable required preload before Catapult can read
      ADDR_WIDTH     : INTEGER RANGE 12 TO 32 := 32;          -- AXI4-Lite host address width
      DATA_WIDTH     : INTEGER RANGE 32 TO 64 := 32           -- AXI4-Lite host data width (must be 32 or 64)
    );
    PORT(
      -- AXI-4 Lite Interface
      ACLK       : IN   std_logic;                                 -- AXI-4 Bus Clock - Rising edge
      ARESETn    : IN   std_logic;                                 -- Active LOW synchronous reset
      -- ============== AXI4-Lite Write Address Channel Signals
      AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);               -- Write address
      AWVALID    : IN   std_logic;                                          -- Write address valid
      AWREADY    : OUT  std_logic;                                          -- Write address ready (slave is ready to accept AWADDR)
      -- ============== AXI4-Lite Write Data Channel
      WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0); -- Write data
      WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise) - ignored in AXI-4 Lite
      WVALID     : IN   std_logic;                                          -- Write data is valid
      WREADY     : OUT  std_logic;                                          -- Write ready (slave is ready to accept WDATA)
      -- ============== AXI4-Lite Write Response Channel Signals
      BRESP      : OUT  std_logic_vector(1 downto 0);                       -- Write response (of slave) - only OKAY, SLVERR, DECERR supported in AXI-4 Lite
      BVALID     : OUT  std_logic;                                          -- Write response valid (slave accepted WDATA)
      BREADY     : IN   std_logic;                                          -- Response ready (master can accept slave's write response)
      -- ============== AXI4-Lite Read Address Channel Signals
      ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);               -- Read address
      ARVALID    : IN   std_logic;                                          -- Read address valid
      ARREADY    : OUT  std_logic;                                          -- Read address ready (slave is ready to accept ARADDR)
      -- ============== AXI4-Lite Read Data Channel Signals
      RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0); -- Read data
      RRESP      : OUT  std_logic_vector(1 downto 0);                       -- Read response (of slave) - only OKAY, SLVERR, DECERR supported in AXI-4 Lite
      RVALID     : OUT  std_logic;                                          -- Read valid (slave providing RDATA)
      RREADY     : IN   std_logic;                                          -- Read ready (master ready to receive RDATA)

      -- Catapult interface assuming sidebyside packing 
      clk        : IN   std_logic;                                     -- Catapult Clock
      arst_n     : IN   std_logic;                                     -- Reset
--    d_from_ccs : IN   std_logic_vector(cwidth-1 downto 0);           -- Data out of Catapult block
--    d_from_vld : IN   std_logic;                                     -- Data out is valid
      d_to_ccs   : OUT  std_logic_vector(cwidth-1 downto 0)            -- Data into Catapult bloc
    );
  END COMPONENT;

  
  -- AXI4 Lite Slave Output
  COMPONENT ccs_axi4_lite_slave_out
    GENERIC(
      rscid          : INTEGER               := 1;            -- Required resource ID parameter
      op_width       : INTEGER RANGE 1 TO 64 := 1;            -- Operator width (dummy parameter)
      cwidth         : INTEGER RANGE 1 TO 256 := 32;          -- Internal register width
      nopreload      : INTEGER RANGE 0 TO 1 := 0;             -- 1=disable required preload before Catapult can read
      ADDR_WIDTH     : INTEGER RANGE 12 TO 32 := 32;          -- AXI4-Lite host address width
      DATA_WIDTH     : INTEGER RANGE 32 TO 64 := 32           -- AXI4-Lite host data width (must be 32 or 64)
    );
    PORT(
      -- AXI-4 Lite Interface
      ACLK       : IN   std_logic;                                     -- AXI-4 Bus Clock - Rising edge
      ARESETn    : IN   std_logic;                                     -- Active LOW synchronous reset
      -- ============== AXI4-Lite Write Address Channel Signals
      AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Write address
      AWVALID    : IN   std_logic;                                     -- Write address valid
      AWREADY    : OUT  std_logic;                                     -- Write address ready (slave is ready to accept AWADDR)
      --AWLEN      : IN   std_logic_vector(7 downto 0);                -- Write burst length    - must always be 0 in AXI4-Lite
      --AWSIZE     : IN   std_logic_vector(1 downto 0);                -- Write burst size      - must equal host_dw_bytes-2
      --AWBURST    : IN   std_logic_vector(1 downto 0);                -- Write burst mode      - must always be 0 (fixed mode) in AXI4-Lite
      --AWLOCK     : IN   std_logic;                                   -- Lock type             - must always be 0 (Normal access) in AXI4-Lite
      --AWCACHE    : IN   std_logic_vector(3 downto 0);                -- Memory type           - must always be 0 (Non-modifiable, Non-bufferable) in AXI4-Lite
      --AWPROT     : IN   std_logic_vector(2 downto 0);                -- Protection Type       - ignored in this model
      -- ============== AXI4-Lite Write Data Channel
      WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);       -- Write data
      WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise) - ignored in AXI-4 Lite
      WVALID     : IN   std_logic;                                     -- Write data is valid
      WREADY     : OUT  std_logic;                                     -- Write ready (slave is ready to accept WDATA)
      -- ============== AXI4-Lite Write Response Channel Signals
      BRESP      : OUT  std_logic_vector(1 downto 0);                  -- Write response (of slave) - only OKAY, SLVERR, DECERR supported in AXI-4 Lite
      BVALID     : OUT  std_logic;                                     -- Write response valid (slave accepted WDATA)
      BREADY     : IN   std_logic;                                     -- Response ready (master can accept slave's write response)
      -- ============== AXI4-Lite Read Address Channel Signals
      ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Read address
      ARVALID    : IN   std_logic;                                     -- Read address valid
      ARREADY    : OUT  std_logic;                                     -- Read address ready (slave is ready to accept ARADDR)
      --ARLEN      : IN   std_logic_vector(7 downto 0);                -- Read burst length     - must always be 0 in AXI4-Lite
      --ARSIZE     : IN   std_logic_vector(1 downto 0);                -- Read burst size       - must equal host_dw_bytes-2
      --ARBURST    : IN   std_logic_vector(1 downto 0);                -- Read burst mode       - must always be 0 (fixed mode) in AXI4-Lite
      --ARLOCK     : IN   std_logic;                                   -- Lock type             - must always be 0 (Normal access) in AXI4-Lite
      --ARCACHE    : IN   std_logic_vector(3 downto 0);                -- Memory type           - must always be 0 (Non-modifiable, Non-bufferable) in AXI4-Lite
      --ARPROT     : IN   std_logic_vector(2 downto 0);                -- Protection Type       - ignored in this model
      -- ============== AXI4-Lite Read Data Channel Signals
      RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);       -- Read data
      RRESP      : OUT  std_logic_vector(1 downto 0);                  -- Read response (of slave) - only OKAY, SLVERR, DECERR supported in AXI-4 Lite
      RVALID     : OUT  std_logic;                                     -- Read valid (slave providing RDATA)
      RREADY     : IN   std_logic;                                     -- Read ready (master ready to receive RDATA)

      -- Catapult interface assuming sidebyside packing 
      d_from_ccs : IN   std_logic_vector(cwidth-1 downto 0);           -- Data out of Catapult block
      d_from_vld : IN   std_logic                                      -- Data out is valid
--    d_to_ccs   : OUT  std_logic_vector(cwidth-1 downto 0)            -- Data into Catapult bloc
    );
  END COMPONENT;

  COMPONENT ccs_axi4_slave_mem
    GENERIC(
      rscid           : integer                 := 1;    -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;   -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;    -- dummy parameter for cwidth calculation
      cwidth          : integer range 1 to 1024 := 8;    -- Internal memory data width
      addr_w          : integer range 1 to 64   := 4;    -- Catapult address bus widths
      nopreload       : integer range 0 to 1    := 0;    -- 1= no preload before Catapult can read
      rst_ph          : integer range 0 to 1    := 0;    -- Reset phase.  1= Positive edge. Default is AXI negative edge
      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;   -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;   -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;    -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;    -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;    -- AXI4 Region Map (ignored in this model)
      wBASE_ADDRESS   : integer                 := 0;    -- AXI4 write channel base address alignment based on data bus width
      rBASE_ADDRESS   : integer                 := 0     -- AXI4 read channel base address alignment based on data bus width
     );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                     -- Rising edge clock
      ARESETn    : IN   std_logic;                                     -- Active LOW asynchronous reset

      -- ============== AXI4 Write Address Channel Signals
      AWID       : IN   std_logic_vector(ID_WIDTH-1 downto 0);         -- Write address ID
      AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Write address
      AWLEN      : IN   std_logic_vector(7 downto 0);                  -- Write burst length
      AWSIZE     : IN   std_logic_vector(2 downto 0);                  -- Write burst size
      AWBURST    : IN   std_logic_vector(1 downto 0);                  -- Write burst mode
      AWLOCK     : IN   std_logic;                                     -- Lock type
      AWCACHE    : IN   std_logic_vector(3 downto 0);                  -- Memory type
      AWPROT     : IN   std_logic_vector(2 downto 0);                  -- Protection Type
      AWQOS      : IN   std_logic_vector(3 downto 0);                  -- Quality of Service
      AWREGION   : IN   std_logic_vector(3 downto 0);                  -- Region identifier
      AWUSER     : IN   std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
      AWVALID    : IN   std_logic;                                     -- Write address valid
      AWREADY    : OUT  std_logic;                                     -- Write address ready (slave is ready to accept AWADDR)

      -- ============== AXI4 Write Data Channel
      WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);       -- Write data
      WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise)
      WLAST      : IN   std_logic;                                     -- Write last
      WUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
      WVALID     : IN   std_logic;                                     -- Write data is valid
      WREADY     : OUT  std_logic;                                     -- Write ready (slave is ready to accept WDATA)
      
      -- ============== AXI4 Write Response Channel Signals
      BID        : OUT  std_logic_vector(ID_WIDTH-1 downto 0);         -- Response ID tag
      BRESP      : OUT  std_logic_vector(1 downto 0);                  -- Write response (of slave)
      BUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
      BVALID     : OUT  std_logic;                                     -- Write response valid (slave accepted WDATA)
      BREADY     : IN   std_logic;                                     -- Response ready (master can accept slave's write response)
      
      -- ============== AXI4 Read Address Channel Signals
      ARID       : IN   std_logic_vector(ID_WIDTH-1 downto 0);         -- Read address ID
      ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Read address
      ARLEN      : IN   std_logic_vector(7 downto 0);                  -- Read burst length
      ARSIZE     : IN   std_logic_vector(2 downto 0);                  -- Read burst size
      ARBURST    : IN   std_logic_vector(1 downto 0);                  -- Read burst mode
      ARLOCK     : IN   std_logic;                                     -- Lock type
      ARCACHE    : IN   std_logic_vector(3 downto 0);                  -- Memory type
      ARPROT     : IN   std_logic_vector(2 downto 0);                  -- Protection Type
      ARQOS      : IN   std_logic_vector(3 downto 0);                  -- Quality of Service
      ARREGION   : IN   std_logic_vector(3 downto 0);                  -- Region identifier
      ARUSER     : IN   std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
      ARVALID    : IN   std_logic;                                     -- Read address valid
      ARREADY    : OUT  std_logic;                                     -- Read address ready (slave is ready to accept ARADDR)
      
      -- ============== AXI4 Read Data Channel Signals
      RID        : OUT  std_logic_vector(ID_WIDTH-1 downto 0);         -- Read ID tag
      RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);       -- Read data
      RRESP      : OUT  std_logic_vector(1 downto 0);                  -- Read response (of slave)
      RLAST      : OUT  std_logic;                                     -- Read last
      RUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
      RVALID     : OUT  std_logic;                                     -- Read valid (slave providing RDATA)
      RREADY     : IN   std_logic;                                     -- Read ready (master ready to receive RDATA)
      
      -- Catapult interface
      s_re      : IN   std_logic;                                      -- Catapult attempting read of slave memory
      s_we      : IN   std_logic;                                      -- Catapult attempting write to slave memory
      s_raddr   : IN   std_logic_vector(addr_w-1 downto 0);            -- Catapult addressing into memory (axi_addr = base_addr + s_raddr)
      s_waddr   : IN   std_logic_vector(addr_w-1 downto 0);            -- Catapult addressing into memory (axi_addr = base_addr + s_waddr)
      s_din     : OUT  std_logic_vector(cwidth-1 downto 0);            -- Data into catapult block through this interface
      s_dout    : IN   std_logic_vector(cwidth-1 downto 0);            -- Data out to slave from catapult
      s_rrdy    : OUT  std_logic;                                      -- Read data is valid
      s_wrdy    : OUT  std_logic;                                      -- Slave memory ready for write by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                      -- component is idle - clock can be suppressed
      tr_write_done : IN std_logic;                                    -- transactor resource preload write done
      s_tdone   : IN   std_logic                                       -- Transaction_done in scverify
    );  
  END COMPONENT;

  COMPONENT ccs_axi4_master_read_core
    GENERIC(
      rscid           : integer                 := 1;      -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;     -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 1 to 64   := 4;      -- Catapult address bus width
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      xburstsize      : integer                 := 0;      -- Burst size for scverify transactor
      xBASE_ADDRESS   : integer                 := 0;      -- Base address for scverify transactor
      xBASE_ADDRESSU  : integer                 := 0       -- Upper word for 64-bit Base address for scverify transactor
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset
      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready
      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- Configuration interface
      cfgBaseAddress : IN  std_logic_vector(ADDR_WIDTH-1 downto 0);  
      cfgBurstSize   : IN  std_logic_vector(31 downto 0);            
      cfgTimeout     : IN  std_logic_vector(31 downto 0);            

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_raddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for read request (axi_addr = base_addr + m_raddr)
      m_rburst  : IN   std_logic_vector(31 downto 0);                   -- Read Burst length (constant rburstsize for now, future enhancement driven by operator)
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic                                        -- The component is idle. The next clk can be suppressed
    );
  END COMPONENT;
  
  COMPONENT ccs_axi4_master_read
    GENERIC(
      rscid           : integer                 := 1;      -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;     -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 1 to 64   := 4;      -- Catapult address bus width
      burstsize       : integer                 := 0;      -- Catapult configuration option for Read burst size
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      timeout         : integer                 := 0;      --  #cycles timeout for burst stall

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      BASE_ADDRESS    : integer                 := 0;      -- Base address 
      BASE_ADDRESSU   : integer                 := 0       -- Upper word for 64-bit Base address 
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset
      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready
      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_raddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for read request (axi_addr = base_addr + m_raddr)
      m_rburst  : IN   std_logic_vector(31 downto 0);                   -- Read Burst length (constant rburstsize for now, future enhancement driven by operator)
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic                                        -- The component is idle. The next clk can be suppressed
    );
  END COMPONENT;
  
  COMPONENT ccs_axi4_master_write_core
    GENERIC(
      rscid           : integer                 := 1;      -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;     -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 1 to 64   := 4;      -- Catapult address bus width
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      xburstsize      : integer                 := 0;      -- Burst size for scverify transactor
      xBASE_ADDRESS   : integer                 := 0;      -- Base address for scverify transactor
      xBASE_ADDRESSU  : integer                 := 0       -- Upper word for 64-bit Base address for scverify transactor
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset

      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);                   -- Write burst length
      AWSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Write burst size
      AWBURST    : OUT  std_logic_vector(1 downto 0);                   -- Write burst mode
      AWLOCK     : OUT  std_logic;                                      -- Lock type
      AWCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      AWPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      AWQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      AWUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      AWVALID    : OUT  std_logic;                                      -- Write address valid
      AWREADY    : IN   std_logic;                                      -- Write address ready

      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);        -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);    -- Write strobe (bytewise)
      WLAST      : OUT  std_logic;                                      -- Write last
      WUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      WVALID     : OUT  std_logic;                                      -- Write data is valid
      WREADY     : IN   std_logic;                                      -- Write ready

      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);                   -- Write response
      BUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      BVALID     : IN   std_logic;                                      -- Write response valid
      BREADY     : OUT  std_logic;                                      -- Response ready

      -- Configuration interface
      cfgBaseAddress : IN  std_logic_vector(ADDR_WIDTH-1 downto 0);  
      cfgBurstSize   : IN  std_logic_vector(31 downto 0);            
      cfgTimeout     : IN  std_logic_vector(31 downto 0);            

      -- Catapult interface
      m_we      : IN   std_logic;                                       -- Catapult attempting write to memory over bus
      m_waddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for write request (axi_addr = base_addr + m_waddr)
      m_wburst  : IN   std_logic_vector(31 downto 0);                   -- Write Burst length (constant wburstsize for now, future enhancement driven by operator)
      m_dout    : IN   std_logic_vector(cwidth-1 downto 0);             -- Data out to bus from catapult (write request)
      m_wrdy    : OUT  std_logic;                                       -- Bus memory ready for write access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      -- Transactor resource interface (for SCVerify simulation only)
      m_wCaughtUp : OUT  std_logic;                                     -- wburst_in == wburst_out
      m_wstate    : OUT  std_logic_vector(2 downto 0)                   -- write_state of master
    );
  END COMPONENT;
  
  COMPONENT ccs_axi4_master_write
    GENERIC(
      rscid           : integer                 := 1;      -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;     -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 1 to 64   := 4;      -- Catapult address bus width
      burstsize       : integer                 := 0;      -- Catapult configuration option for write burst size
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      timeout         : integer                 := 0;      --  #cycles timeout for burst stall

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      BASE_ADDRESS    : integer                 := 0;      -- Base address
      BASE_ADDRESSU   : integer                 := 0       -- Upper word for 64-bit Base address
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset

      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);                   -- Write burst length
      AWSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Write burst size
      AWBURST    : OUT  std_logic_vector(1 downto 0);                   -- Write burst mode
      AWLOCK     : OUT  std_logic;                                      -- Lock type
      AWCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      AWPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      AWQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      AWUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      AWVALID    : OUT  std_logic;                                      -- Write address valid
      AWREADY    : IN   std_logic;                                      -- Write address ready

      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);        -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);    -- Write strobe (bytewise)
      WLAST      : OUT  std_logic;                                      -- Write last
      WUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      WVALID     : OUT  std_logic;                                      -- Write data is valid
      WREADY     : IN   std_logic;                                      -- Write ready

      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);                   -- Write response
      BUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      BVALID     : IN   std_logic;                                      -- Write response valid
      BREADY     : OUT  std_logic;                                      -- Response ready

      -- Catapult interface
      m_we      : IN   std_logic;                                       -- Catapult attempting write to memory over bus
      m_waddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for write request (axi_addr = base_addr + m_waddr)
      m_wburst  : IN   std_logic_vector(31 downto 0);                   -- Write Burst length (constant wburstsize for now, future enhancement driven by operator)
      m_dout    : IN   std_logic_vector(cwidth-1 downto 0);             -- Data out to bus from catapult (write request)
      m_wrdy    : OUT  std_logic;                                       -- Bus memory ready for write access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      -- Transactor resource interface (for SCVerify simulation only)
      m_wCaughtUp : OUT  std_logic;                                     -- wburst_in == wburst_out
      m_wstate    : OUT  std_logic_vector(2 downto 0)                   -- write_state of master
    );
  END COMPONENT;
  
  COMPONENT ccs_axi4_master_core
    GENERIC(
      rscid           : integer                 := 1;      -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;     -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 1 to 64   := 4;      -- Catapult address bus width
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      xwburstsize     : integer                 := 0;      -- wBurst size for scverify transactor
      xrburstsize     : integer                 := 0;      -- rBurst size for scverify transactor
      xwBASE_ADDRESS  : integer                 := 0;      -- wBase address for scverify transactor
      xrBASE_ADDRESS  : integer                 := 0;      -- rBase address for scverify transactor
      xwBASE_ADDRESSU : integer                 := 0;      -- Upper word for 64-bit wBase address for scverify transactor
      xrBASE_ADDRESSU : integer                 := 0       -- Upper word for 64-bit rBase address for scverify transactor
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset
      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);                   -- Write burst length
      AWSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Write burst size
      AWBURST    : OUT  std_logic_vector(1 downto 0);                   -- Write burst mode
      AWLOCK     : OUT  std_logic;                                      -- Lock type
      AWCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      AWPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      AWQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      AWUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      AWVALID    : OUT  std_logic;                                      -- Write address valid
      AWREADY    : IN   std_logic;                                      -- Write address ready
      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);        -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);    -- Write strobe (bytewise)
      WLAST      : OUT  std_logic;                                      -- Write last
      WUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      WVALID     : OUT  std_logic;                                      -- Write data is valid
      WREADY     : IN   std_logic;                                      -- Write ready
      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);                   -- Write response
      BUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      BVALID     : IN   std_logic;                                      -- Write response valid
      BREADY     : OUT  std_logic;                                      -- Response ready
      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready
      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- Configuration interface
      cfgwBaseAddress : IN  std_logic_vector(ADDR_WIDTH-1 downto 0);  
      cfgrBaseAddress : IN  std_logic_vector(ADDR_WIDTH-1 downto 0);  
      cfgwBurstSize  : IN  std_logic_vector(31 downto 0);            
      cfgrBurstSize  : IN  std_logic_vector(31 downto 0);            
      cfgTimeout     : IN  std_logic_vector(31 downto 0);

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_we      : IN   std_logic;                                       -- Catapult attempting write to memory over bus
      m_waddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for write request (axi_addr = base_addr + m_waddr)
      m_raddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for read request (axi_addr = base_addr + m_raddr)
      m_wburst  : IN   std_logic_vector(31 downto 0);                   -- Write Burst length (constant wburstsize for now, future enhancement driven by operator)
      m_rburst  : IN   std_logic_vector(31 downto 0);                   -- Read Burst length (constant rburstsize for now, future enhancement driven by operator)
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_dout    : IN   std_logic_vector(cwidth-1 downto 0);             -- Data out to bus from catapult (write request)
      m_wrdy    : OUT  std_logic;                                       -- Bus memory ready for write access by Catapult (1=ready)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      -- Transactor resource interface (for SCVerify simulation only)
      m_wCaughtUp : OUT  std_logic;                                     -- wburst_in == wburst_out
      m_wstate    : OUT  std_logic_vector(2 downto 0)                   -- write_state of master
    );
  END COMPONENT;

  COMPONENT ccs_axi4_master_cfg
    GENERIC(
      rscid           : integer                 := 1;      -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;     -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 1 to 64   := 4;      -- Catapult address bus width
      cburst_mode     : integer range 0 to 2    := 0;      -- Burst mode (0==use w/rburstsize, 1==configuration port)
      wburstsize      : integer                 := 0;      -- Catapult configuration option for Write burst size
      rburstsize      : integer                 := 0;      -- Catapult configuration option for Read burst size
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      use_go          : integer range 0 to 1    := 0;      -- Use the cfgBus stop/go mechanism.  Default not.

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      base_addr_mode  : integer range 0 to 2    := 0;      -- Where base address is specified (0=param, 1=cfg, 2=port)
      wBASE_ADDRESS   : integer                 := 0;      -- AXI4 write channel base address
      rBASE_ADDRESS   : integer                 := 0;      -- AXI4 read channel base address
      wBASE_ADDRESSU  : integer                 := 0;      -- Upper word of 64-bit AXI4 write channel base address
      rBASE_ADDRESSU  : integer                 := 0       -- Upper word of 64-bit AXI4 read channel base address
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset
      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);                   -- Write burst length
      AWSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Write burst size
      AWBURST    : OUT  std_logic_vector(1 downto 0);                   -- Write burst mode
      AWLOCK     : OUT  std_logic;                                      -- Lock type
      AWCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      AWPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      AWQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      AWUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      AWVALID    : OUT  std_logic;                                      -- Write address valid
      AWREADY    : IN   std_logic;                                      -- Write address ready
      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);        -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);    -- Write strobe (bytewise)
      WLAST      : OUT  std_logic;                                      -- Write last
      WUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      WVALID     : OUT  std_logic;                                      -- Write data is valid
      WREADY     : IN   std_logic;                                      -- Write ready
      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);                   -- Write response
      BUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      BVALID     : IN   std_logic;                                      -- Write response valid
      BREADY     : OUT  std_logic;                                      -- Response ready
      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready
      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- AXI-lite slave interface to program base_addr - address 0, 1, 2
      cfgAWADDR  : IN  std_logic_vector(31 downto 0);
      cfgAWVALID : IN  std_logic;
      cfgAWREADY : OUT std_logic;
      cfgWDATA   : IN  std_logic_vector(31 downto 0);
      cfgWSTRB   : IN  std_logic_vector(3 downto 0);
      cfgWVALID  : IN  std_logic;
      cfgWREADY  : OUT std_logic;
      cfgBRESP   : OUT std_logic_vector(1 downto 0);
      cfgBVALID  : OUT std_logic;
      cfgBREADY  : IN  std_logic;
      cfgARADDR  : IN  std_logic_vector(31 downto 0);
      cfgARVALID : IN  std_logic;
      cfgARREADY : OUT std_logic;
      cfgRDATA   : OUT std_logic_vector(31 downto 0);
      cfgRRESP   : OUT std_logic_vector(1 downto 0);
      cfgRVALID  : OUT std_logic;
      cfgRREADY  : IN  std_logic;

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_we      : IN   std_logic;                                       -- Catapult attempting write to memory over bus
      m_waddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for write request (axi_addr = base_addr + m_waddr)
      m_raddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for read request (axi_addr = base_addr + m_raddr)
      m_wburst  : IN   std_logic_vector(31 downto 0);                   -- Write Burst length (constant wburstsize for now, future enhancement driven by operator)
      m_rburst  : IN   std_logic_vector(31 downto 0);                   -- Read Burst length (constant rburstsize for now, future enhancement driven by operator)
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_dout    : IN   std_logic_vector(cwidth-1 downto 0);             -- Data out to bus from catapult (write request)
      m_wrdy    : OUT  std_logic;                                       -- Bus memory ready for write access by Catapult (1=ready)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      -- Transactor resource interface (for SCVerify simulation only)
      m_wCaughtUp : OUT  std_logic;                                     -- wburst_in == wburst_out
      m_wstate    : OUT  std_logic_vector(2 downto 0)                   -- write_state of master
    );
  END COMPONENT;

  COMPONENT ccs_axi4_master
    GENERIC(
      rscid           : integer                 := 1;      -- Resource ID
      -- Catapult Bus Configuration generics
      depth           : integer                 := 16;     -- Number of addressable elements (up to 20bit address)
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 1 to 64   := 4;      -- Catapult address bus width
      wburstsize      : integer                 := 0;      -- Catapult configuration option for Write burst size
      rburstsize      : integer                 := 0;      -- Catapult configuration option for Read burst size
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      timeout         : integer                 := 0;      --  #cycles timeout for burst stall

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      wBASE_ADDRESS    : integer                := 0;      -- AXI4 write channel base address
      rBASE_ADDRESS    : integer                := 0;      -- AXI4 read channel base address
      wBASE_ADDRESSU   : integer                := 0;      -- Upper word for 64-bit AXI4 write channel base address
      rBASE_ADDRESSU   : integer                := 0       -- Upper word for 64-bit AXI4 read channel base addressable
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset
      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);                   -- Write burst length
      AWSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Write burst size
      AWBURST    : OUT  std_logic_vector(1 downto 0);                   -- Write burst mode
      AWLOCK     : OUT  std_logic;                                      -- Lock type
      AWCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      AWPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      AWQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      AWUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      AWVALID    : OUT  std_logic;                                      -- Write address valid
      AWREADY    : IN   std_logic;                                      -- Write address ready
      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);        -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);    -- Write strobe (bytewise)
      WLAST      : OUT  std_logic;                                      -- Write last
      WUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      WVALID     : OUT  std_logic;                                      -- Write data is valid
      WREADY     : IN   std_logic;                                      -- Write ready
      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);                   -- Write response
      BUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      BVALID     : IN   std_logic;                                      -- Write response valid
      BREADY     : OUT  std_logic;                                      -- Response ready
      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready
      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_we      : IN   std_logic;                                       -- Catapult attempting write to memory over bus
      m_waddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for write request (axi_addr = base_addr + m_waddr)
      m_raddr   : IN   std_logic_vector(addr_w    -1 downto 0);         -- Address for read request (axi_addr = base_addr + m_raddr)
      m_wburst  : IN   std_logic_vector(31 downto 0);                   -- Write Burst length (constant wburstsize for now, future enhancement driven by operator)
      m_rburst  : IN   std_logic_vector(31 downto 0);                   -- Read Burst length (constant rburstsize for now, future enhancement driven by operator)
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_dout    : IN   std_logic_vector(cwidth-1 downto 0);             -- Data out to bus from catapult (write request)
      m_wrdy    : OUT  std_logic;                                       -- Bus memory ready for write access by Catapult (1=ready)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      -- Transactor resource interface (for SCVerify simulation only)
      m_wCaughtUp : OUT  std_logic;                                     -- wburst_in == wburst_out
      m_wstate    : OUT  std_logic_vector(2 downto 0)                   -- write_state of master
    );
  END COMPONENT;

COMPONENT ccs_axi4_master_instream_core
    GENERIC(
      rscid           : integer                 := 1;     -- Resource ID
      -- Catapult Bus Configuration generics
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 0 to 64   := 4;      -- Catapult address bus width
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      fpga            : integer range 0 to 1    := 0;      -- Choose the fpga better-route version
      
      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      xburstsize      : integer                 := 0;      -- Burst size for scverify transactor
      xframe_size      : integer                := 16;     -- Number of elements in the frame to be streamed
      xBASE_ADDRESS   : integer                 := 0;      -- Base address for scverify transactor
      xBASE_ADDRESSU  : integer                 := 0       -- Upper word for 64-bit Base address for scverify transactor
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset

      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready

      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- Configuration interface
      cfgBaseAddress : IN  std_logic_vector(ADDR_WIDTH-1 downto 0);  
      cfgBurstSize   : IN  std_logic_vector(31 downto 0);            
      cfgTimeout     : IN  std_logic_vector(31 downto 0);            
      cfgFrameSize   : IN  std_logic_vector(31 downto 0);            

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      rdy       : OUT  std_logic                                        -- For transactor
    );

END COMPONENT;

COMPONENT ccs_axi4_master_outstream_core
    GENERIC(
      rscid           : integer;                           -- Resource ID
      -- Catapult Bus Configuration generics
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 0 to 64   := 4;      -- Catapult address bus width
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16   := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      xburstsize       : integer                := 0;      -- Burst size for scverify transactor
      xframe_size      : integer                := 16;     -- Number of elements in the frame to be streamed
      xBASE_ADDRESS    : integer                := 0;      -- Base addess  for scverify transactor
      xBASE_ADDRESSU   : integer                := 0       -- Upper word for 64-bit Base addess  for scverify transactor
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset

      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);                   -- Write burst length
      AWSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Write burst size
      AWBURST    : OUT  std_logic_vector(1 downto 0);                   -- Write burst mode
      AWLOCK     : OUT  std_logic;                                      -- Lock type
      AWCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      AWPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      AWQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      AWUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      AWVALID    : OUT  std_logic;                                      -- Write address valid
      AWREADY    : IN   std_logic;                                      -- Write address ready

      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);        -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);    -- Write strobe (bytewise)
      WLAST      : OUT  std_logic;                                      -- Write last
      WUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      WVALID     : OUT  std_logic;                                      -- Write data is valid
      WREADY     : IN   std_logic;                                      -- Write ready

      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);                   -- Write response
      BUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      BVALID     : IN   std_logic;                                      -- Write response valid
      BREADY     : OUT  std_logic;                                      -- Response ready

      -- Catapult interface
      -- Configuration interface
      cfgBaseAddress : IN  std_logic_vector(ADDR_WIDTH-1 downto 0);  
      cfgBurstSize   : IN  std_logic_vector(31 downto 0);            
      cfgTimeout     : IN  std_logic_vector(31 downto 0);            
      cfgFrameSize   : IN  std_logic_vector(31 downto 0);            

      m_we      : IN   std_logic;                                       -- Catapult attempting write to memory over bus
      m_dout    : IN   std_logic_vector(cwidth-1 downto 0);             -- Data out to bus from catapult (write request)
      m_wrdy    : OUT  std_logic;                                       -- Bus memory ready for write access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      vld       : OUT  std_logic                                        -- Core produced data.  Written into transactor "row"
    );

END COMPONENT;

COMPONENT ccs_axi4_master_instream
    GENERIC(
      rscid           : integer                 := 1;     -- Resource ID
      -- Catapult Bus Configuration generics
      frame_size      : integer                 := 16;     -- Number of elements in the frame to be streamed
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 0 to 64   := 4;      -- Catapult address bus width
      burstsize       : integer                 := 0;      -- Catapult configuration option for Read burst size
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      fpga            : integer range 0 to 1    := 0;      -- Choose the fpga better-route version
      timeout         : integer                 := 0;      --  #cycles timeout for burst stall
      
      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      BASE_ADDRESS    : integer                 := 0;      -- Base address 
      BASE_ADDRESSU   : integer                 := 0       -- Upper word for 64-bit Base address 
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset

      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready

      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      rdy       : OUT  std_logic                                        -- For transactor
    );

END COMPONENT;

COMPONENT ccs_axi4_master_outstream
    GENERIC(
      rscid           : integer;                           -- Resource ID
      -- Catapult Bus Configuration generics
      frame_size      : integer                 := 16;     -- Number of elements in the frame to be streamed
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 0 to 64   := 4;      -- Catapult address bus width
      burstsize       : integer                 := 0;      -- Catapult configuration option for Write burst size
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      timeout         : integer                 := 0;      --  #cycles timeout for burst stall

      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16   := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;     -- AXI4 Region Map (ignored in this model)
      BASE_ADDRESS    : integer                := 0;      -- AXI4 write channel base address
      BASE_ADDRESSU   : integer                := 0       -- Upper word for 64-bit AXI4 write channel base address
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset

      -- ============== AXI4 Write Address Channel Signals
      AWID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Write address ID
      AWADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Write address
      AWLEN      : OUT  std_logic_vector(7 downto 0);                   -- Write burst length
      AWSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Write burst size
      AWBURST    : OUT  std_logic_vector(1 downto 0);                   -- Write burst mode
      AWLOCK     : OUT  std_logic;                                      -- Lock type
      AWCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      AWPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      AWQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      AWREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      AWUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      AWVALID    : OUT  std_logic;                                      -- Write address valid
      AWREADY    : IN   std_logic;                                      -- Write address ready

      -- ============== AXI4 Write Data Channel
      WDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);        -- Write data
      WSTRB      : OUT  std_logic_vector((DATA_WIDTH/8)-1 downto 0);    -- Write strobe (bytewise)
      WLAST      : OUT  std_logic;                                      -- Write last
      WUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      WVALID     : OUT  std_logic;                                      -- Write data is valid
      WREADY     : IN   std_logic;                                      -- Write ready

      -- ============== AXI4 Write Response Channel Signals
      BID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Response ID tag
      BRESP      : IN   std_logic_vector(1 downto 0);                   -- Write response
      BUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      BVALID     : IN   std_logic;                                      -- Write response valid
      BREADY     : OUT  std_logic;                                      -- Response ready

      -- Catapult interface
      m_we      : IN   std_logic;                                       -- Catapult attempting write to memory over bus
      m_dout    : IN   std_logic_vector(cwidth-1 downto 0);             -- Data out to bus from catapult (write request)
      m_wrdy    : OUT  std_logic;                                       -- Bus memory ready for write access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      vld       : OUT  std_logic                                        -- Core produced data.  Written into transactor "row"
    );

END COMPONENT;

COMPONENT ccs_axi4_lite_slave_outreg
  GENERIC(
    rscid           : integer                 := 1;    -- Resource ID
    -- Catapult Bus Configuration generics
    op_width        : integer range 1 to 1024 := 1;    -- dummy parameter for cwidth calculation
    cwidth          : integer range 1 to 1024 := 8;    -- Internal memory data width
    rst_ph          : integer range 0 to 1    := 0;    -- Reset phase.  1= Positive edge. Default is AXI negative edge
    -- AXI-4 Bus Configuration generics
    ADDR_WIDTH      : integer range 12 to 64  := 32;   -- AXI4 bus address width
    DATA_WIDTH      : integer range 8 to 1024 := 32;   -- AXI4 read&write data bus width
    BASE_ADDRESS   : integer                  := 0     -- AXI4 Address that the register is seen at
    );
  PORT(
    -- AXI-4 Interface
    ACLK       : IN   std_logic;                                     -- Rising edge clock
    ARESETn    : IN   std_logic;                                     -- Active LOW asynchronous reset
    
    -- ============== AXI4 Read Address Channel Signals
    ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Read address
    ARVALID    : IN   std_logic;                                     -- Read address valid
    ARREADY    : OUT  std_logic;                                     -- Read address ready (slave is ready to accept ARADDR)
    
    -- ============== AXI4 Read Data Channel Signals
    RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);       -- Read data
    RRESP      : OUT  std_logic_vector(1 downto 0);                  -- Read response (of slave)
    RVALID     : OUT  std_logic;                                     -- Read valid (slave providing RDATA)
    RREADY     : IN   std_logic;                                     -- Read ready (master ready to receive RDATA)
    
    -- Catapult interface
    ivld      : IN   std_logic;                                      -- Catapult data ready
    idat      : in   std_logic_vector(cwidth-1 downto 0);            -- Data from catapult

    -- External valid flag
    vld       : OUT  std_logic                                       -- Data valid for AXI read
    );

END COMPONENT;

COMPONENT ccs_axi4_lite_slave_inreg 
  GENERIC(
    rscid           : integer                 := 1;    -- Resource ID
    -- Catapult Bus Configuration generics
    op_width        : integer range 1 to 1024 := 1;    -- dummy parameter for cwidth calculation
    cwidth          : integer range 1 to 1024 := 8;    -- Internal memory data width
    rst_ph          : integer range 0 to 1    := 0;    -- Reset phase.  1= Positive edge. Default is AXI negative edge
    disable_vld     : integer range 0 to 1    := 0;    -- Disable use of vld signal to stall I/O
    -- AXI-4 Bus Configuration generics
    ADDR_WIDTH      : integer range 12 to 64  := 32;   -- AXI4 bus address width
    DATA_WIDTH      : integer range 8 to 1024 := 32;   -- AXI4 read&write data bus width
    BASE_ADDRESS    : integer                 := 0     -- AXI4 Address that the register is seen at
    );
  PORT(
    -- AXI-4 Interface
    ACLK       : IN   std_logic;                                     -- Rising edge clock
    ARESETn    : IN   std_logic;                                     -- Active LOW asynchronous reset
    -- ============== AXI4 Write Address Channel Signals
    AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Write address
    AWVALID    : IN   std_logic;                                     -- Write address valid
    AWREADY    : OUT  std_logic;                                     -- Write address ready (slave is ready to accept AWADDR)
    -- ============== AXI4 Write Data Channel
    WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);       -- Write data
    WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise)
    WVALID     : IN   std_logic;                                     -- Write data is valid
    WREADY     : OUT  std_logic;                                     -- Write ready (slave is ready to accept WDATA)
    
    -- ============== AXI4 Write Response Channel Signals
    BRESP      : OUT  std_logic_vector(1 downto 0);                  -- Write response (of slave)
    BVALID     : OUT  std_logic;                                     -- Write response valid (slave accepted WDATA)
    BREADY     : IN   std_logic;                                     -- Response ready (master can accept slave's write response)
    
    -- Catapult interface
    ivld      : OUT   std_logic;                                      -- Data valid.  Duration 1 cycle
    idat      : OUT   std_logic_vector(cwidth-1 downto 0)             -- Data into catapult block through this interface
    );
END COMPONENT;

COMPONENT ccs_axi4_lite_slave_indirect
  GENERIC(
    rscid           : integer                 := 1;    -- Resource ID
    -- Catapult Bus Configuration generics
    op_width        : integer range 1 to 1024 := 1;    -- dummy parameter for cwidth calculation
    cwidth          : integer range 1 to 1024 := 8;    -- Internal memory data width
    rst_ph          : integer range 0 to 1    := 0;    -- Reset phase.  1= Positive edge. Default is AXI negative edge
    -- AXI-4 Bus Configuration generics
    ADDR_WIDTH      : integer range 12 to 64  := 32;   -- AXI4 bus address width
    DATA_WIDTH      : integer range 8 to 1024 := 32;   -- AXI4 read&write data bus width
    BASE_ADDRESS    : integer                 := 0     -- AXI4 Address that the register is seen at
    );
  PORT(
    -- AXI-4 Interface
    ACLK       : IN   std_logic;                                     -- Rising edge clock
    ARESETn    : IN   std_logic;                                     -- Active LOW asynchronous reset
    -- ============== AXI4 Write Address Channel Signals
    AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Write address
    AWVALID    : IN   std_logic;                                     -- Write address valid
    AWREADY    : OUT  std_logic;                                     -- Write address ready (slave is ready to accept AWADDR)
    -- ============== AXI4 Write Data Channel
    WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);       -- Write data
    WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise)
    WVALID     : IN   std_logic;                                     -- Write data is valid
    WREADY     : OUT  std_logic;                                     -- Write ready (slave is ready to accept WDATA)
    
    -- ============== AXI4 Write Response Channel Signals
    BRESP      : OUT  std_logic_vector(1 downto 0);                  -- Write response (of slave)
    BVALID     : OUT  std_logic;                                     -- Write response valid (slave accepted WDATA)
    BREADY     : IN   std_logic;                                     -- Response ready (master can accept slave's write response)
    
    -- ============== AXI4 Read Address Channel Signals
    ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Read address
    ARVALID    : IN   std_logic;                                     -- Read address valid
    ARREADY    : OUT  std_logic;                                     -- Read address ready (slave is ready to accept ARADDR)
    
    -- ============== AXI4 Read Data Channel Signals
    RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);       -- Read data
    RRESP      : OUT  std_logic_vector(1 downto 0);                  -- Read response (of slave)
    RVALID     : OUT  std_logic;                                     -- Read valid (slave providing RDATA)
    RREADY     : IN   std_logic;                                     -- Read ready (master ready to receive RDATA)
    
    -- Catapult interface
    idat      : OUT   std_logic_vector(cwidth-1 downto 0)             -- Data into catapult block through this interface
    );
END COMPONENT;

COMPONENT ccs_axi4_lite_slave_outsync
  GENERIC(
    rscid           : integer                 := 1;    -- Resource ID
    -- Catapult Bus Configuration generics
    rst_ph          : integer range 0 to 1    := 0;    -- Reset phase.  1= Positive edge. Default is AXI negative edge
    -- AXI-4 Bus Configuration generics
    ADDR_WIDTH      : integer range 12 to 32  := 32;   -- AXI4 bus address width
    DATA_WIDTH      : integer range 32 to 64  := 32;   -- AXI4 read&write data bus width
    BASE_ADDRESS   : integer                  := 0     -- AXI4 Address that the register is seen at
    );
  PORT(
    -- AXI-4 Interface
    ACLK       : IN   std_logic;                                     -- Rising edge clock
    ARESETn    : IN   std_logic;                                     -- Active LOW asynchronous reset
    
    -- ============== AXI4 Write Address Channel Signals
    AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Write address
    AWVALID    : IN   std_logic;                                     -- Write address valid
    AWREADY    : OUT  std_logic;                                     -- Write address ready (slave is ready to accept AWADDR)

    -- ============== AXI4 Write Data Channel
    WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);       -- Write data
    WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe - not used in LITE
    WVALID     : IN   std_logic;                                     -- Write data is valid
    WREADY     : OUT  std_logic;                                     -- Write ready (slave is ready to accept WDATA)
    
    -- ============== AXI4 Write Response Channel Signals
    BRESP      : OUT  std_logic_vector(1 downto 0);                  -- Write response (of slave)
    BVALID     : OUT  std_logic;                                     -- Write response valid (slave accepted WDATA)
    BREADY     : IN   std_logic;                                     -- Response ready (master can accept slave's write response)
    
    -- ============== AXI4 Read Address Channel Signals
    ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Read address
    ARVALID    : IN   std_logic;                                     -- Read address valid
    ARREADY    : OUT  std_logic;                                     -- Read address ready (slave is ready to accept ARADDR)
    
    -- ============== AXI4 Read Data Channel Signals
    RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);       -- Read data
    RRESP      : OUT  std_logic_vector(1 downto 0);                  -- Read response (of slave)
    RVALID     : OUT  std_logic;                                     -- Read valid (slave providing RDATA)
    RREADY     : IN   std_logic;                                     -- Read ready (master ready to receive RDATA)
    
    -- Catapult interface
    irdy      : OUT  std_logic;                                      -- Catapult data ready
    ivld      : IN   std_logic;                                      -- Catapult data ready
    triosy    : OUT  std_logic                                       -- Data from catapult
    );

END COMPONENT;

COMPONENT ccs_axi4_lite_slave_insync
  GENERIC(
    rscid           : integer                 := 1;    -- Resource ID
    -- Catapult Bus Configuration generics
    rst_ph          : integer range 0 to 1    := 0;    -- Reset phase.  1= Positive edge. Default is AXI negative edge
    -- AXI-4 Bus Configuration generics
    ADDR_WIDTH      : integer range 12 to 32  := 32;   -- AXI4 bus address width
    DATA_WIDTH      : integer range 32 to 64  := 32;   -- AXI4 read&write data bus width
    BASE_ADDRESS    : integer                 := 0     -- AXI4 Address that the register is seen at
    );
  PORT(
    -- AXI-4 Interface
    ACLK       : IN   std_logic;                                     -- Rising edge clock
    ARESETn    : IN   std_logic;                                     -- Active LOW asynchronous reset
    -- ============== AXI4 Write Address Channel Signals
    AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Write address
    AWVALID    : IN   std_logic;                                     -- Write address valid
    AWREADY    : OUT  std_logic;                                     -- Write address ready (slave is ready to accept AWADDR)
    -- ============== AXI4 Write Data Channel
    WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);       -- Write data
    WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise)
    WVALID     : IN   std_logic;                                     -- Write data is valid
    WREADY     : OUT  std_logic;                                     -- Write ready (slave is ready to accept WDATA)
    
    -- ============== AXI4 Write Response Channel Signals
    BRESP      : OUT  std_logic_vector(1 downto 0);                  -- Write response (of slave)
    BVALID     : OUT  std_logic;                                     -- Write response valid (slave accepted WDATA)
    BREADY     : IN   std_logic;                                     -- Response ready (master can accept slave's write response)
    
    -- ============== AXI4 Read Address Channel Signals
    ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Read address
    ARVALID    : IN   std_logic;                                     -- Read address valid
    ARREADY    : OUT  std_logic;                                     -- Read address ready (slave is ready to accept ARADDR)
    
    -- ============== AXI4 Read Data Channel Signals
    RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);       -- Read data
    RRESP      : OUT  std_logic_vector(1 downto 0);                  -- Read response (of slave)
    RVALID     : OUT  std_logic;                                     -- Read valid (slave providing RDATA)
    RREADY     : IN   std_logic;                                     -- Read ready (master ready to receive RDATA)

    -- Catapult interface
    irdy      : IN    std_logic;
    ivld      : OUT   std_logic;
    triosy    : OUT   std_logic                                       -- // transactor uses 
    );
END COMPONENT;


  -- ==============================================================
  -- APB Components

  -- Used to define the APB bus definition (direction of signals is from the slave's perspective)
  COMPONENT apb_busdef
    GENERIC(
      width        : INTEGER RANGE 1 TO 32 := 32;           -- Number of bits in an element
      addr_width   : INTEGER RANGE 1 TO 32 := 1             -- Number of address bits to address 'words' elements
    );
    PORT(
      -- APB interface
      PCLK      : IN   std_logic;                           -- Rising edge clock
      PRESETn   : IN   std_logic;                           -- Active LOW synchronous reset
      PADDR     : IN   std_logic_vector(addr_width-1 downto 0);  -- APB Bridge driven address bus (32 bit max)
      PSELx     : IN   std_logic;                           -- APB Bridge driven select for this slave
      PWRITE    : IN   std_logic;                           -- APB Bridge driven read/write signal (0=read)
      PENABLE   : IN   std_logic;                           -- APB Bridge driven enable signal
      PWDATA    : IN   std_logic_vector(width-1 downto 0);  -- APB Bridge driven data to write to slave (32 bit max)
      PRDATA    : OUT  std_logic_vector(width-1 downto 0);  -- Slave driven data back to APB Bridge (32 bit max)
      PREADY    : OUT  std_logic;                           -- Slave driven signal to extend transfer cycles (1=ready)
      PSLVERR   : OUT  std_logic                            -- Slave driven signal indicating transfer failed (1=fail)
    );
  END COMPONENT;

  COMPONENT apb_master
    GENERIC(
      words        : INTEGER RANGE 1 TO 256 := 1;           -- Number of addressable elements
      width        : INTEGER RANGE 1 TO 32 := 32;           -- Number of bits in an element
      addr_width   : INTEGER RANGE 1 TO 32 := 1             -- Number of address bits to address 'words' elements
    );
    PORT(
      -- APB interface
      PCLK      : IN   std_logic;                           -- Rising edge clock
      PRESETn   : IN   std_logic;                           -- Active LOW synchronous reset
      PADDR     : OUT  std_logic_vector(30 downto 0);       -- APB Bridge driven address bus (32 bit max)
      PSELx     : OUT  std_logic;                           -- APB Bridge driven select for this slave
      PWRITE    : OUT  std_logic;                           -- APB Bridge driven read/write signal (0=read)
      PENABLE   : OUT  std_logic;                           -- APB Bridge driven enable signal
      PWDATA    : OUT  std_logic_vector(width-1 downto 0);  -- APB Bridge driven data to write to slave (32 bit max)
      PRDATA    : IN   std_logic_vector(width-1 downto 0);  -- Slave driven data back to APB Bridge (32 bit max)
      PREADY    : IN   std_logic;                           -- Slave driven signal to extend transfer cycles (1=ready)
      PSLVERR   : IN   std_logic;                           -- Slave driven signal indicating transfer failed (1=fail)
      -- Catapult interface
      m_rw      : IN   std_logic;                           -- read/write
      m_strobe  : IN   std_logic;                           -- initiate a bus transfer
      m_adr     : IN   std_logic_vector(addr_width-1 downto 0); -- target address
      m_din     : OUT  std_logic_vector(width-1 downto 0);  -- data in from slave
      m_dout    : IN   std_logic_vector(width-1 downto 0);  -- data out to slave
      m_rdy     : OUT  std_logic                            -- ready for transfer (1=ready)
    );
  END COMPONENT;

  -- APB slave memory
  COMPONENT apb_slave_mem
    GENERIC(
      words          : INTEGER RANGE 1 TO 256 := 1;            -- Number of addressable elements
      width          : INTEGER RANGE 1 TO 32 := 32;           -- Number of bits in an element
      addr_width     : INTEGER RANGE 1 TO 32 := 1;            -- Number of address bits to address 'words' elements
      num_rwports    : INTEGER RANGE 1 TO 100 := 1;           -- Number of register file "ports"
      nopreload      : INTEGER RANGE 0 TO 1 := 0              -- 1=disable required preload before Catapult can read
    );
    PORT(
      -- APB interface
      PCLK      : IN   std_logic;                           -- Rising edge clock
      PRESETn   : IN   std_logic;                           -- Active LOW synchronous reset
      PADDR     : IN   std_logic_vector(30 downto 0);       -- APB Bridge driven address bus (32 bit max)
      PSELx     : IN   std_logic;                           -- APB Bridge driven select for this slave
      PWRITE    : IN   std_logic;                           -- APB Bridge driven read/write signal (0=read)
      PENABLE   : IN   std_logic;                           -- APB Bridge driven enable signal
      PWDATA    : IN   std_logic_vector(width-1 downto 0);  -- APB Bridge driven data to write to slave (32 bit max)
      PRDATA    : OUT  std_logic_vector(width-1 downto 0);  -- Slave driven data back to APB Bridge (32 bit max)
      PREADY    : OUT  std_logic;                           -- Slave driven signal to extend transfer cycles (1=ready)
      PSLVERR   : OUT  std_logic;                           -- Slave driven signal indicating transfer failed (1=fail)
      -- Catapult interface
      s_rw      : IN   std_logic_vector(num_rwports-1 downto 0);            -- read/write
      s_strobe  : IN   std_logic_vector(num_rwports-1 downto 0);            -- Catapult attempting read of slave
      s_adr     : IN   std_logic_vector(num_rwports*addr_width-1 downto 0); -- Catapult addressing into memory
      s_din     : OUT  std_logic_vector(num_rwports*width-1 downto 0);      -- Data into catapult block through this interface
      s_dout    : IN   std_logic_vector(num_rwports*width-1 downto 0);      -- Data out to slave from catapult
      s_rdy     : OUT  std_logic_vector(num_rwports-1 downto 0)             -- Slave memory ready for read (1=ready)
    );
  END COMPONENT;

  -- ==============================================================
  -- Internally referenced components

  COMPONENT amba_generic_reg
    GENERIC (
      width    : INTEGER := 1;
      ph_en    : INTEGER RANGE 0 TO 1 := 1;
      has_en   : INTEGER RANGE 0 TO 1 := 1
    );
    PORT (
      clk     : IN  std_logic;
      en      : IN  std_logic;
      arst    : IN  std_logic;
      srst    : IN  std_logic;
      d       : IN  std_logic_vector(width-1 DOWNTO 0);
      z       : OUT std_logic_vector(width-1 DOWNTO 0)
    );
  END COMPONENT;

  COMPONENT amba_pipe_ctrl
    GENERIC (
      rscid    : INTEGER := 0;
      width    : INTEGER := 8;
      sz_width : INTEGER := 8;
      fifo_sz  : INTEGER RANGE 0 TO 128 := 8;
      ph_en    : INTEGER RANGE 0 TO 1 := 1
    );
    PORT (
      clk      : IN  std_logic;
      en       : IN  std_logic;
      arst     : IN  std_logic;
      srst     : IN  std_logic;
      din_vld  : IN  std_logic;
      din_rdy  : OUT std_logic;
      din      : IN  std_logic_vector(width-1 DOWNTO 0);
      dout_vld : OUT std_logic;
      dout_rdy : IN  std_logic;
      dout     : OUT std_logic_vector(width-1 DOWNTO 0);
      sd       : OUT std_logic_vector(sz_width-1 DOWNTO 0)
    );
  END COMPONENT;

  COMPONENT amba_pipe
    GENERIC (
      rscid    : INTEGER := 0;
      width    : INTEGER := 8;
      sz_width : INTEGER := 8;
      fifo_sz  : INTEGER RANGE 0 TO 128 := 8;
      ph_en    : INTEGER RANGE 0 TO 1 := 1
    );
    PORT (
      -- clock
      clk      : IN  std_logic;
      en       : IN  std_logic;
      arst     : IN  std_logic;
      srst     : IN  std_logic;
      -- writer
      din_rdy  : OUT std_logic;
      din_vld  : IN  std_logic;
      din      : IN  std_logic_vector(width-1 DOWNTO 0);
      -- reader
      dout_rdy : IN  std_logic;
      dout_vld : OUT std_logic;
      dout     : OUT std_logic_vector(width-1 DOWNTO 0);
      -- size
      sz       : OUT std_logic_vector(sz_width-1 DOWNTO 0);
      sz_req   : in  std_logic
    );
  END COMPONENT;

  COMPONENT amba_ctrl_in_buf_wait
    GENERIC (
      width    : INTEGER := 8
    );
    PORT (
      clk      : IN  std_logic;
      arst     : IN  std_logic;
      irdy   : IN  std_logic;
      ivld   : OUT std_logic;
      idat   : OUT std_logic_vector(width-1 DOWNTO 0);
      rdy    : OUT std_logic;
      vld    : IN  std_logic;
      dat    : IN  std_logic_vector(width-1 DOWNTO 0);
      is_idle : out std_logic
    );
  END COMPONENT;

  COMPONENT ML_amba_ctrl_in_buf_wait
    GENERIC (
      width    : INTEGER := 8
    );
    PORT (
      clk      : IN  std_logic;
      arst     : IN  std_logic;
      irdy   : IN  std_logic;
      ivld   : OUT std_logic;
      idat   : OUT std_logic_vector(width-1 DOWNTO 0);
      rdy    : OUT std_logic;
      vld    : IN  std_logic;
      dat    : IN  std_logic_vector(width-1 DOWNTO 0);
      is_idle : out std_logic
    );
  END COMPONENT;

COMPONENT ML_ccs_axi4_master_fpga_instream_core
    GENERIC(
      rscid           : integer                 := 1;     -- Resource ID
      -- Catapult Bus Configuration generics
      frame_size      : integer                 := 16;     -- Number of elements in the frame to be streamed
      op_width        : integer range 1 to 1024 := 1;      -- dummy parameter for cwidth calculation
      cwidth          : integer range 8 to 1024 := 32;     -- Catapult data bus width (multiples of 8)
      addr_w          : integer range 0 to 64   := 4;      -- Catapult address bus width
      rst_ph          : integer range 0 to 1    := 0;      -- Reset phase - negative default
      
      -- AXI-4 Bus Configuration generics
      ADDR_WIDTH      : integer range 12 to 64  := 32;     -- AXI4 bus address width
      DATA_WIDTH      : integer range 8 to 1024 := 32;     -- AXI4 read&write data bus width
      ID_WIDTH        : integer range 1 to 16    := 1;      -- AXI4 ID field width (ignored in this model)
      USER_WIDTH      : integer range 1 to 32   := 1;      -- AXI4 User field width (ignored in this model)
      REGION_MAP_SIZE : integer range 1 to 15   := 1;      -- AXI4 Region Map (ignored in this model)
      xburstsize      : integer                 := 0;      -- Burst size for scverify transactor
      xBASE_ADDRESS   : integer                 := 0;      -- Base address for scverify transactor
      xBASE_ADDRESSU  : integer                 := 0       -- Upper word for 64-bit Base address for scverify transactor
    );
    PORT(
      -- AXI-4 Interface
      ACLK       : IN   std_logic;                                      -- Rising edge clock
      ARESETn    : IN   std_logic;                                      -- Active LOW asynchronous reset

      -- ============== AXI4 Read Address Channel Signals
      ARID       : OUT  std_logic_vector(ID_WIDTH-1 downto 0);          -- Read address ID
      ARADDR     : OUT  std_logic_vector(ADDR_WIDTH-1 downto 0);        -- Read address
      ARLEN      : OUT  std_logic_vector(7 downto 0);                   -- Read burst length
      ARSIZE     : OUT  std_logic_vector(2 downto 0);                   -- Read burst size
      ARBURST    : OUT  std_logic_vector(1 downto 0);                   -- Read burst mode
      ARLOCK     : OUT  std_logic;                                      -- Lock type
      ARCACHE    : OUT  std_logic_vector(3 downto 0);                   -- Memory type
      ARPROT     : OUT  std_logic_vector(2 downto 0);                   -- Protection Type
      ARQOS      : OUT  std_logic_vector(3 downto 0);                   -- Quality of Service
      ARREGION   : OUT  std_logic_vector(3 downto 0);                   -- Region identifier
      ARUSER     : OUT  std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      ARVALID    : OUT  std_logic;                                      -- Read address valid
      ARREADY    : IN   std_logic;                                      -- Read address ready

      -- ============== AXI4 Read Data Channel Signals
      RID        : IN   std_logic_vector(ID_WIDTH-1 downto 0);          -- Read ID tag
      RDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);        -- Read data
      RRESP      : IN   std_logic_vector(1 downto 0);                   -- Read response
      RLAST      : IN   std_logic;                                      -- Read last
      RUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);        -- User signal
      RVALID     : IN   std_logic;                                      -- Read valid
      RREADY     : OUT  std_logic;                                      -- Read ready

      -- Configuration interface
      cfgBaseAddress : IN  std_logic_vector(ADDR_WIDTH-1 downto 0);  
      cfgBurstSize   : IN  std_logic_vector(31 downto 0);            
      cfgTimeout     : IN  std_logic_vector(31 downto 0);            

      -- Catapult interface
      m_re      : IN   std_logic;                                       -- Catapult attempting read of memory over bus
      m_din     : OUT  std_logic_vector(cwidth-1 downto 0);             -- Data into catapult block through this interface (read request)
      m_rrdy    : OUT  std_logic;                                       -- Bus memory ready for read access by Catapult (1=ready)
      is_idle   : OUT  std_logic;                                       -- The component is idle. The next clk can be suppressed
      rdy       : OUT  std_logic                                        -- For transactor
    );
END COMPONENT;

  
  -- ==============================================================
  -- AMBA Protocol Constants

  -- AxBURST modes
  CONSTANT AXI4_AxBURST_FIXED    : std_logic_vector(1 downto 0) := "00";
  CONSTANT AXI4_AxBURST_INCR     : std_logic_vector(1 downto 0) := "01";
  CONSTANT AXI4_AxBURST_WRAP     : std_logic_vector(1 downto 0) := "10";
  CONSTANT AXI4_AxBURST_RESERVED : std_logic_vector(1 downto 0) := "11";
  -- AxLOCK modes
  CONSTANT AXI4_AxLOCK_NORMAL    : std_logic                    := '0';
  CONSTANT AXI4_AxLOCK_EXCLUSIVE : std_logic                    := '1';
  -- Memory types W and R mostly the xame
  CONSTANT AXI4_AWCACHE_NB        : std_logic_vector(3 downto 0) := "0000";
  CONSTANT AXI4_AWCACHE_B         : std_logic_vector(3 downto 0) := "0001";
  CONSTANT AXI4_AWCACHE_NORM_NCNB : std_logic_vector(3 downto 0) := "0010"; --
  CONSTANT AXI4_AWCACHE_NORM_NCB  : std_logic_vector(3 downto 0) := "0011" ;
  CONSTANT AXI4_AWCACHE_WTNA      : std_logic_vector(3 downto 0) := "0110";
  CONSTANT AXI4_AWCACHE_WTRA      : std_logic_vector(3 downto 0) := "0110";
  CONSTANT AXI4_AWCACHE_WTWA      : std_logic_vector(3 downto 0) := "1110";
  CONSTANT AXI4_AWCACHE_WTRWA     : std_logic_vector(3 downto 0) := "1110";
  CONSTANT AXI4_AWCACHE_WBNA      : std_logic_vector(3 downto 0) := "0111";
  CONSTANT AXI4_AWCACHE_WBRA      : std_logic_vector(3 downto 0) := "0111";
  CONSTANT AXI4_WACACHE_WBWA      : std_logic_vector(3 downto 0) := "1111";
  CONSTANT AXI4_AWCACHE_WBRWA     : std_logic_vector(3 downto 0) := "1111";
  CONSTANT AXI4_ARCACHE_NB        : std_logic_vector(3 downto 0) := "0000";
  CONSTANT AXI4_ARCACHE_B         : std_logic_vector(3 downto 0) := "0001";
  CONSTANT AXI4_ARCACHE_NORM_NCNB : std_logic_vector(3 downto 0) := "0010"; --
  CONSTANT AXI4_ARCACHE_NORM_NCB  : std_logic_vector(3 downto 0) := "0011" ;
  CONSTANT AXI4_ARCACHE_WTNA      : std_logic_vector(3 downto 0) := "1010";
  CONSTANT AXI4_ARCACHE_WTRA      : std_logic_vector(3 downto 0) := "1110";
  CONSTANT AXI4_ARCACHE_WTWA      : std_logic_vector(3 downto 0) := "1010";
  CONSTANT AXI4_ARCACHE_WTRWA     : std_logic_vector(3 downto 0) := "1110";
  CONSTANT AXI4_ARCACHE_WBNA      : std_logic_vector(3 downto 0) := "1011";
  CONSTANT AXI4_ARCACHE_WBRA      : std_logic_vector(3 downto 0) := "1111";
  CONSTANT AXI4_ARCACHE_WBWA      : std_logic_vector(3 downto 0) := "1011";
  CONSTANT AXI4_ARCACHE_WBRWA     : std_logic_vector(3 downto 0) := "1111";
  -- QOS pre-defines
  CONSTANT AXI4_AxQOS_NONE        : std_logic_vector(3 downto 0) := "0000";
  -- AxSIZE byte sizes
  CONSTANT AXI4_AxSIZE_001_BYTE  : std_logic_vector(2 downto 0) := "000";
  CONSTANT AXI4_AxSIZE_002_BYTE  : std_logic_vector(2 downto 0) := "001";
  CONSTANT AXI4_AxSIZE_004_BYTE  : std_logic_vector(2 downto 0) := "010";
  CONSTANT AXI4_AxSIZE_008_BYTE  : std_logic_vector(2 downto 0) := "011";
  CONSTANT AXI4_AxSIZE_016_BYTE  : std_logic_vector(2 downto 0) := "100";
  CONSTANT AXI4_AxSIZE_032_BYTE  : std_logic_vector(2 downto 0) := "101";
  CONSTANT AXI4_AxSIZE_064_BYTE  : std_logic_vector(2 downto 0) := "110";
  CONSTANT AXI4_AxSIZE_128_BYTE  : std_logic_vector(2 downto 0) := "111";
  -- AxPROT bit fields
  CONSTANT AXI4_AxPROT_b0_UNPRIV   : std_logic := '0';
  CONSTANT AXI4_AxPROT_b0_PRIV     : std_logic := '1';
  CONSTANT AXI4_AxPROT_b1_SECURE   : std_logic := '0';
  CONSTANT AXI4_AxPROT_b1_UNSECURE : std_logic := '1';
  CONSTANT AXI4_AxPROT_b2_DATA     : std_logic := '0';
  CONSTANT AXI4_AxPROT_b2_INSTR    : std_logic := '1';
  -- xRESP response codes
  CONSTANT AXI4_xRESP_OKAY         : std_logic_vector(1 downto 0) := "00";
  CONSTANT AXI4_xRESP_EXOKAY       : std_logic_vector(1 downto 0) := "01";
  CONSTANT AXI4_xRESP_SLVERR       : std_logic_vector(1 downto 0) := "10";
  CONSTANT AXI4_xRESP_DECERR       : std_logic_vector(1 downto 0) := "11";

  -- Utility function(s) to support debug needs
  FUNCTION bits ( size : INTEGER) RETURN INTEGER;
  FUNCTION slv2bin(vec: std_logic_vector) RETURN string;
  FUNCTION slv2hex(vec: std_logic_vector) RETURN string;

END PACKAGE amba_comps;

PACKAGE BODY amba_comps IS

   -- Find the number of bits required to represent an unsigned
   -- number less than size
  FUNCTION bits (size : integer) RETURN INTEGER IS
  BEGIN
    IF (size < 0) THEN RETURN 0;
    ELSIF (size = 0) THEN RETURN 1;
    ELSE
      FOR i IN 1 TO size LOOP
        IF (2**i >= size) THEN
          RETURN i;
        END IF;
      END LOOP;
      RETURN 0;
    END IF;
  END;

   -- Convert an std_logic_vector to a (hex)string for printing
   -- vec needs to be a multiple of 4 in size
  FUNCTION slv2hex(vec: std_logic_vector) RETURN string IS
      variable quad : std_logic_vector(3 downto 0);
      constant ne: integer := vec'length/4;
      variable s: string(1 to ne);
   BEGIN
      if vec'length mod 4 /= 0 then
         assert false
         report "slv2hex called with slv lenght that is not a multiple of 4";
         return s;
      end if;
      for i in 0 to ne-1 loop
         quad := vec(4*i+3 downto 4*i);
         case quad is
            when x"0" => s(ne-i) := '0';
            when x"1" => s(ne-i) := '1';
            when x"2" => s(ne-i) := '2';
            when x"3" => s(ne-i) := '3';
            when x"4" => s(ne-i) := '4';
            when x"5" => s(ne-i) := '5';
            when x"6" => s(ne-i) := '6';
            when x"7" => s(ne-i) := '7';
            when x"8" => s(ne-i) := '8';
            when x"9" => s(ne-i) := '9';
            when x"A" => s(ne-i) := 'A';
            when x"B" => s(ne-i) := 'B';
            when x"C" => s(ne-i) := 'C';
            when x"D" => s(ne-i) := 'D';
            when x"E" => s(ne-i) := 'E';
            when x"F" => s(ne-i) := 'F';
            when others => s(ne-i) := '-';
         end case;
      end loop;
      return s;
   END;

   -- Convert an std_logic_vector to a (binary)string for printing
   FUNCTION slv2bin(vec: std_logic_vector) RETURN string IS
      VARIABLE stmp: string(vec'left+1 downto 1);
   BEGIN
      FOR i in vec'reverse_range LOOP
         IF (vec(i) = 'U') THEN
            stmp(i+1) := 'U';
         ELSIF (vec(i) = 'X') THEN
            stmp(i+1) := 'X';
         ELSIF (vec(i) = '0') THEN
            stmp(i+1) := '0';
         ELSIF (vec(i) = '1') THEN
            stmp(i+1) := '1';
         ELSIF (vec(i) = 'Z') THEN
            stmp(i+1) := 'Z';
         ELSIF (vec(i) = 'W') THEN
            stmp(i+1) := 'W';
         ELSIF (vec(i) = 'L') THEN
            stmp(i+1) := 'L';
         ELSIF (vec(i) = 'H') THEN
            stmp(i+1) := 'H';
         ELSE
            stmp(i+1) := '-';
         END IF;
      END LOOP;
      RETURN stmp;
   END;

END amba_comps;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/ccs_libs/interfaces/amba/ccs_axi4_slave_mem.vhd 

-- --------------------------------------------------------------------------
-- DESIGN UNIT:        ccs_axi4_slave_mem
--
-- DESCRIPTION:
--   This model implements an AXI-4 Slave memory interface for use in 
--   Interface Synthesis in Catapult. The component details are described in the datasheet.
--
--   AXI/Catapult read/write to the same address in the same cycle is non-determinant
--
-- Notes:
--  1. This model implements a local memory of size {cwidth x depth}.
--     If the Catapult operation requires a memory width cwidth <= AXI bus width
--     this model will zero-pad the high end bits as necessary.
-- CHANGE LOG:
--  01/29/19 - Add reset phase and separate base address for read/write channels
--  11/26/18 - Add burst and other tweaks
--  02/28/18 - Initial implementation
--
-- -------------------------------------------------------------------------------
--  Memory Organization
--   This model is designed to provide storage for only the bits/elements that
--   the Catapult core actually interacts with.
--   The user supplies a base address for the AXI memory store via BASE_ADDRESS
--   parameter.  
-- Example:
--   C++ array declared as "ac_int<7,false>  coeffs[4];"
--   results in a Catapult operator width (op_width) of 7,
--   and cwidth=7 and addr_w=2 (addressing 4 element locations).
--   The library forces DATA_WIDTH to be big enough to hold
--   cwidth bits, rounded up to power-of-2 as needed.
--
--   The AXI address scheme addresses bytes and so increments
--   by number-of-bytes per data transaction, plus the BASE_ADDRESS. 
--   The top and left describe the AXI view of the memory. 
--   The bottom and right describe the Catapult view of the memory.
--
--      AXI-4 SIGNALS
--      ADDR_WIDTH=4        DATA_WIDTH=32
--        AxADDR               xDATA
--                    31                       0
--                    +------------+-----------+
--      BA+0000       |            |           |
--                    +------------+-----------+
--      BA+0000       |            |           |
--                    +------------+===========+
--      BA+1100       |            |  elem3    |    11
--                    +------------+===========+
--      BA+1000       |            |  elem2    |    10
--                    +------------+===========+
--      BA+0100       |            |  elem1    |    01
--                    +------------+===========+
--      BA+0000       |            |  elem0    |    00
--                    +------------+===========+
--                                 6           0
--                                   s_din/out     s_addr
--                                   cwidth=7      addr_w=2
--                                         CATAPULT SIGNALS
--
-- -------------------------------------------------------------------------------

LIBRARY ieee;

  USE ieee.std_logic_1164.all;
  USE ieee.numeric_std.all;       
  USE std.textio.all;
  USE ieee.std_logic_textio.all;
  USE ieee.math_real.all;


USE work.amba_comps.all;

ENTITY ccs_axi4_slave_mem IS
  GENERIC(
    rscid           : integer                 := 1;    -- Resource ID
    -- Catapult Bus Configuration generics
    depth           : integer                 := 16;   -- Number of addressable elements (up to 20bit address)
    op_width        : integer range 1 to 1024 := 1;    -- dummy parameter for cwidth calculation
    cwidth          : integer range 1 to 1024 := 8;    -- Internal memory data width
    addr_w          : integer range 1 to 64   := 4;    -- Catapult address bus widths
    nopreload       : integer range 0 to 1    := 0;    -- 1= no preload before Catapult can read
    rst_ph          : integer range 0 to 1    := 0;    -- Reset phase.  1= Positive edge. Default is AXI negative edge
    -- AXI-4 Bus Configuration generics
    ADDR_WIDTH      : integer range 12 to 64  := 32;   -- AXI4 bus address width
    DATA_WIDTH      : integer range 8 to 1024 := 32;   -- AXI4 read&write data bus width
    ID_WIDTH        : integer range 1 to 16   := 1;    -- AXI4 ID field width (ignored in this model)
    USER_WIDTH      : integer range 1 to 32   := 1;    -- AXI4 User field width (ignored in this model)
    REGION_MAP_SIZE : integer range 1 to 15   := 1;    -- AXI4 Region Map (ignored in this model)
    wBASE_ADDRESS   : integer                 := 0;    -- AXI4 write channel base address alignment based on data bus width
    rBASE_ADDRESS   : integer                 := 0     -- AXI4 read channel base address alignment based on data bus width
    );
  PORT(
    -- AXI-4 Interface
    ACLK       : IN   std_logic;                                     -- Rising edge clock
    ARESETn    : IN   std_logic;                                     -- Active LOW asynchronous reset
    -- ============== AXI4 Write Address Channel Signals
    AWID       : IN   std_logic_vector(ID_WIDTH-1 downto 0);         -- Write address ID
    AWADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Write address
    AWLEN      : IN   std_logic_vector(7 downto 0);                  -- Write burst length
    AWSIZE     : IN   std_logic_vector(2 downto 0);                  -- Write burst size
    AWBURST    : IN   std_logic_vector(1 downto 0);                  -- Write burst mode
    AWLOCK     : IN   std_logic;                                     -- Lock type
    AWCACHE    : IN   std_logic_vector(3 downto 0);                  -- Memory type
    AWPROT     : IN   std_logic_vector(2 downto 0);                  -- Protection Type
    AWQOS      : IN   std_logic_vector(3 downto 0);                  -- Quality of Service
    AWREGION   : IN   std_logic_vector(3 downto 0);                  -- Region identifier
    AWUSER     : IN   std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
    AWVALID    : IN   std_logic;                                     -- Write address valid
    AWREADY    : OUT  std_logic;                                     -- Write address ready (slave is ready to accept AWADDR)
    -- ============== AXI4 Write Data Channel
    WDATA      : IN   std_logic_vector(DATA_WIDTH-1 downto 0);       -- Write data
    WSTRB      : IN   std_logic_vector((DATA_WIDTH/8)-1 downto 0);   -- Write strobe (bytewise)
    WLAST      : IN   std_logic;                                     -- Write last
    WUSER      : IN   std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
    WVALID     : IN   std_logic;                                     -- Write data is valid
    WREADY     : OUT  std_logic;                                     -- Write ready (slave is ready to accept WDATA)
    
    -- ============== AXI4 Write Response Channel Signals
    BID        : OUT  std_logic_vector(ID_WIDTH-1 downto 0);         -- Response ID tag
    BRESP      : OUT  std_logic_vector(1 downto 0);                  -- Write response (of slave)
    BUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
    BVALID     : OUT  std_logic;                                     -- Write response valid (slave accepted WDATA)
    BREADY     : IN   std_logic;                                     -- Response ready (master can accept slave's write response)
    
    -- ============== AXI4 Read Address Channel Signals
    ARID       : IN   std_logic_vector(ID_WIDTH-1 downto 0);         -- Read address ID
    ARADDR     : IN   std_logic_vector(ADDR_WIDTH-1 downto 0);       -- Read address
    ARLEN      : IN   std_logic_vector(7 downto 0);                  -- Read burst length
    ARSIZE     : IN   std_logic_vector(2 downto 0);                  -- Read burst size
    ARBURST    : IN   std_logic_vector(1 downto 0);                  -- Read burst mode
    ARLOCK     : IN   std_logic;                                     -- Lock type
    ARCACHE    : IN   std_logic_vector(3 downto 0);                  -- Memory type
    ARPROT     : IN   std_logic_vector(2 downto 0);                  -- Protection Type
    ARQOS      : IN   std_logic_vector(3 downto 0);                  -- Quality of Service
    ARREGION   : IN   std_logic_vector(3 downto 0);                  -- Region identifier
    ARUSER     : IN   std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
    ARVALID    : IN   std_logic;                                     -- Read address valid
    ARREADY    : OUT  std_logic;                                     -- Read address ready (slave is ready to accept ARADDR)
    
    -- ============== AXI4 Read Data Channel Signals
    RID        : OUT  std_logic_vector(ID_WIDTH-1 downto 0);         -- Read ID tag
    RDATA      : OUT  std_logic_vector(DATA_WIDTH-1 downto 0);       -- Read data
    RRESP      : OUT  std_logic_vector(1 downto 0);                  -- Read response (of slave)
    RLAST      : OUT  std_logic;                                     -- Read last
    RUSER      : OUT  std_logic_vector(USER_WIDTH-1 downto 0);       -- User signal
    RVALID     : OUT  std_logic;                                     -- Read valid (slave providing RDATA)
    RREADY     : IN   std_logic;                                     -- Read ready (master ready to receive RDATA)
    
    -- Catapult interface
    s_re      : IN   std_logic;                                      -- Catapult attempting read of slave memory
    s_we      : IN   std_logic;                                      -- Catapult attempting write to slave memory
    s_raddr   : IN   std_logic_vector(addr_w-1 downto 0);            -- Catapult addressing into memory (axi_addr = base_addr + s_raddr)
    s_waddr   : IN   std_logic_vector(addr_w-1 downto 0);            -- Catapult addressing into memory (axi_addr = base_addr + s_waddr)
    s_din     : OUT  std_logic_vector(cwidth-1 downto 0);            -- Data into catapult block through this interface
    s_dout    : IN   std_logic_vector(cwidth-1 downto 0);            -- Data out to slave from catapult
    s_rrdy    : OUT  std_logic;                                      -- Read data is valid
    s_wrdy    : OUT  std_logic;                                      -- Slave memory ready for write by Catapult (1=ready)
    is_idle   : OUT  std_logic;                                      -- component is idle - clock can be suppressed
    -- Transactor/scverify support
    tr_write_done : IN std_logic;                                    -- transactor resource preload write done
    s_tdone       : IN std_logic                                     -- Transaction_done in scverify
    );
  

    -- Always rule for checking component parameter values
    --  addr_w == bits(depth)
    --    used to ensure that the width of the address bus on the Catapult side
    --    is capable of addressing 'depth' number of elements. 'depth' will be
    --    determined by the array size operator parameter 'size'
    --    (see the PROP_MAP_size attribute)
    --  ADDR_WIDTH >= addr_w
    --    used to ensure that the address width of the Catapult side is
    --    large enough to accommodate the address width of the AXI-4 bus.
    --    (may need some work to align byte addresses)
    --  ADDR_WIDTH >= 32
    --    ensure that the minimum address space is 4k (AXI requirement)
    --  cwidth == 8 + (op_width>8)*8 + (op_width>16)*16 + (op_width>32)*32 + 
    --                (op_width>64)*64 + (op_width>128)*128 + (op_width>256)*256 +
    --                (op_width>512)*512
    --    used to "round up" the operator width 'op_width' to the next power
    --    of two value (8, 16, 32, 64, 128, 256, 512, 1024)
    --    (see the PROP_MAP_width attribute)
    --  DATA_WIDTH >= cwidth
    --    used to ensure that the Catapult data width is large enough to
    --    accommodate the data width of the AXI-4 bus.
    --    - must be power-of-2 bytes.
    --    - #bits must be some positive integer number of bytes.
    --     Note: user can override DATA_WIDTH from the MAP_TO_MODULE
    --     directive during interface synthesis. No checking is done
    --     to ensure that the override value is a power-of-2 bytes.

END ccs_axi4_slave_mem;

ARCHITECTURE rtl of ccs_axi4_slave_mem IS

  -- Signals for current and next state values
  TYPE   read_state_t IS (axi4r_idle, axi4r_read);
  TYPE   write_state_t IS (axi4w_idle, axi4w_write, axi4w_write_done,  axi4w_catwrite, axi4w_catwrite_done);
  SIGNAL read_state       : read_state_t;
  SIGNAL write_state      : write_state_t;

  -- Memory embedded in this slave
  TYPE   mem_type IS ARRAY (depth-1 downto 0) of std_logic_vector(cwidth-1 downto 0);
  SIGNAL mem                : mem_type;


  -- In/out connections and constant outputs  
  SIGNAL AWREADY_reg : std_logic;
  SIGNAL AWID_reg    : std_logic_vector(ID_WIDTH-1 downto 0);
  SIGNAL WREADY_reg  : std_logic;
  SIGNAL BRESP_reg   : std_logic_vector(1 downto 0);
  SIGNAL BVALID_reg  : std_logic;
  SIGNAL ARREADY_reg : std_logic;
  SIGNAL ARID_reg    : std_logic_vector(ID_WIDTH-1 downto 0);
  SIGNAL RDATA_reg   : std_logic_vector(DATA_WIDTH-1 downto 0);
  SIGNAL RRESP_reg   : std_logic_vector(1 downto 0);
  SIGNAL RLAST_reg   : std_logic;
  SIGNAL RVALID_reg  : std_logic;
  SIGNAL s_din_reg   : std_logic_vector(cwidth-1 downto 0);
  SIGNAL s_rrdy_reg  : std_logic;
  SIGNAL s_wrdy_reg  : std_logic;

  SIGNAL rCatOutOfOrder : std_logic;
  SIGNAL catIsReading   : std_logic;
  SIGNAL next_raddr     : integer;
  
  SIGNAL readBurstCnt: std_logic_vector(7 downto 0);   -- how many are left
  SIGNAL wbase_addr   : std_logic_vector(ADDR_WIDTH-1 downto 0);
  SIGNAL rbase_addr   : std_logic_vector(ADDR_WIDTH-1 downto 0);
  SIGNAL address     : std_logic_vector(ADDR_WIDTH-1 downto 0);
  SIGNAL addrShift : integer;
  SIGNAL readAddr : integer;
  SIGNAL writeAddr : integer;
  SIGNAL int_ARESETn : std_logic;
  
-- catapult address sizes are smaller and cause problems used with axi address sizes
  function extCatAddr(catAddr : std_logic_vector(addr_w -1 downto 0))
    return std_logic_vector is
  
    variable axiAddr : std_logic_vector(ADDR_WIDTH-1 downto 0);
  
  begin
    axiAddr := (others => '0');
    axiAddr(addr_w -1 downto 0) := catAddr;
    return axiAddr;
  end function extCatAddr;

BEGIN
  
  int_ARESETn <= ARESETn when (rst_ph = 0) else (not ARESETn);

  addrShift <= 0 when (DATA_WIDTH/8 <= 1)   else 
               1 when (DATA_WIDTH/8 <= 2)   else
               2 when (DATA_WIDTH/8 <= 4)   else
               3 when (DATA_WIDTH/8 <= 8)   else
               4 when (DATA_WIDTH/8 <= 16)  else
               5 when (DATA_WIDTH/8 <= 32)  else
               6 when (DATA_WIDTH/8 <= 64)  else
               7 when (DATA_WIDTH/8 <= 128) else
               0;

  -- unused outputs
  BUSER   <= (others => '0');
  RUSER   <= (others => '0');
  is_idle <= '0';
  
  AWREADY <= AWREADY_reg;
  WREADY  <= WREADY_reg ;
  BID     <= AWID_reg;
  BRESP   <= BRESP_reg  ;
  BVALID  <= BVALID_reg ;
  ARREADY <= ARREADY_reg;
  RID     <= ARID_reg;
  RDATA   <= RDATA_reg  ;
  RRESP   <= RRESP_reg  ;
  RLAST   <= RLAST_reg  ;
  RVALID  <= RVALID_reg ;
  s_din   <= s_din_reg  ;
  s_wrdy  <= s_wrdy_reg and (not s_tdone);
  s_rrdy  <= s_rrdy_reg and (not rCatOutOfOrder);

  wbase_addr <= std_logic_vector(to_unsigned(wBASE_ADDRESS, wbase_addr'length));
  rbase_addr <= std_logic_vector(to_unsigned(rBASE_ADDRESS, rbase_addr'length));
  
  -- pragma translate_off
  -- error checks.  Keep consistent with axi4_master.v/vhd
  -- all data widths the same
  errChk: process
    variable nBytes : std_logic_vector(31 downto 0);
    variable nBytes2 : std_logic_vector(31 downto 0);
  begin  -- process errChk
    nBytes := std_logic_vector(to_unsigned(DATA_WIDTH/8, 32));
    if (cwidth > DATA_WIDTH) then
      report  "Catapult(cwidth=" & integer'image(cwidth) & ") cannot be greater than AXI(DATA_BUS="
        & integer'image(DATA_WIDTH) & ")."
        severity error;
    end if;
    if ( (DATA_WIDTH mod 8) /= 0) then
      report  "Data bus width(DATA_WIDTH=" & integer'image(DATA_WIDTH) & ") not a discrete number of bytes."
        severity error;
    end if;
    if (to_integer(unsigned(nBytes)) = 0) then 
      report  "Data bus width(DATA_WIDTH=" & integer'image(DATA_WIDTH) & ") must be at least 1 byte."
        severity error;
    end if;
    nBytes2 := std_logic_vector(to_unsigned((DATA_WIDTH/8) - 1, 32));
    nBytes2 := nBytes  and nBytes2;
    if ( to_integer(unsigned(nBytes2)) /= 0) then
      report  "Data bus width must be power-of-2 number of bytes(DATA_WIDTH/8=" & integer'image(DATA_WIDTH/8) & ")"
        severity error;
    end if;
    if (ADDR_WIDTH < 12) then
      report  "AXI bus address width(ADDR_WIDTH=" & integer'image(ADDR_WIDTH) & ") must be at least 12 to address 4K memory space."
        severity error;
    end if;
    wait;
  end process errChk;
  -- pragma translate_on
  
  -- AXI4 Bus Read processing
  axiRead: process(ACLK, int_ARESETn)
    -- pragma translate_off
    variable buf : line;
    -- pragma translate_on
    variable useAddr : std_logic_vector(ADDR_WIDTH-1 downto 0);
    variable useAddr2 : std_logic_vector(ADDR_WIDTH-1 downto 0);
  begin
    if (int_ARESETn = '0') then
      read_state <= axi4r_idle;
      ARREADY_reg <= '1';
      ARID_reg <= (others => '0');
      RDATA_reg <= (others => '0');
      RRESP_reg <= AXI4_xRESP_OKAY;
      RLAST_reg <= '0';
      RVALID_reg <= '0';
      readAddr <= 0;
      readBurstCnt <= (others => '0');
    elsif rising_edge(ACLK) then
      if ((read_state = axi4r_idle) and (ARVALID = '1')) then
        useAddr := std_logic_vector(shift_right(unsigned(ARADDR) - unsigned(rbase_addr), addrShift));
        -- Protect from out of range addressing
        if (unsigned(useAddr) < depth) then
          if (cwidth < DATA_WIDTH) then
            RDATA_reg(DATA_WIDTH-1 downto cwidth) <= (others => '0');
            RDATA_reg(cwidth-1 downto 0) <= mem(to_integer(unsigned(useAddr)));
          else
            RDATA_reg <= mem(to_integer(unsigned(useAddr)));
          end if;
          --write(buf, string'("Slave AXI1 read:mem[0x"));
          --write(buf,  slv2hex(useAddr));
          --write(buf, string'("]=0x"));
          --write(buf,  slv2hex(mem(to_integer(unsigned(useAddr)))));
          --write(buf, string'(" at T="));
          --write(buf, now);
          --writeline(output, buf);
        else
          -- pragma translate_off
          write(buf, string'("Error:  Out-of-range AXI memory read access:0x"));
          write(buf,  slv2hex(ARADDR));
          write(buf, string'(" at T="));
          write(buf, now);
          writeline(output, buf);
          -- pragma translate_on
        end if;
        RRESP_reg <= AXI4_xRESP_OKAY;
        readAddr <= to_integer(unsigned(useAddr));
        readBurstCnt <= ARLEN;
        if (unsigned(ARLEN) = 0) then
          ARREADY_reg <= '0';
          RLAST_reg <= '1';
        end if;
        RVALID_reg <= '1';
        ARID_reg <= ARID;
        read_state <= axi4r_read;
      elsif (read_state = axi4r_read) then
        if (RREADY = '1') then
          if (unsigned(readBurstCnt) = 0) then
            -- we already sent the last data
            ARREADY_reg <= '1';
            RRESP_reg <= AXI4_xRESP_OKAY;
            RLAST_reg <= '0';
            RVALID_reg <= '0';
            read_state <= axi4r_idle;               
          else
            useAddr2 := std_logic_vector(to_unsigned(readAddr + 1, useAddr2'length));
            readAddr <= readAddr + 1;
            -- Protect from out of range addressing
            if (unsigned(useAddr2) < depth) then
              if (cwidth < DATA_WIDTH) then
                RDATA_reg(DATA_WIDTH-1 downto cwidth) <= (others => '0');
                RDATA_reg(cwidth-1 downto 0) <=  mem(to_integer(unsigned(useAddr2)));
              else
                RDATA_reg <=  mem(to_integer(unsigned(useAddr2)));
              end if;
              --write(buf, string'("Slave AXI2 read:mem[0x"));
              --write(buf,  slv2hex(useAddr2));
              --write(buf, string'("]=0x"));
              --write(buf,  slv2hex(mem(to_integer(unsigned(useAddr2)))));
              --write(buf, string'(" at T="));
              --write(buf, now);
              --writeline(output, buf);
            else
              -- We bursted right off the end of the array
              -- pragma translate_off
              write(buf, string'("Error:  Out-of-range AXI memory read access:0x"));
              write(buf,  slv2hex(ARADDR));
              write(buf, string'(" at T="));
              write(buf, now);
              writeline(output, buf);
              -- pragma translate_on
            end if;
            readBurstCnt <= std_logic_vector(unsigned(readBurstCnt) - 1);
            if ((unsigned(readBurstCnt) - 1) = 0) then
              ARREADY_reg <= '0';        
              RRESP_reg <= AXI4_xRESP_OKAY;
              RLAST_reg <= '1';
            end if;
            RVALID_reg <= '1';
          end if;
        end if;
      end if;
    end if;
  end process;  -- axiRead process

   -- AXI and catapult write processing.
   -- Catapult write is one-cycle long so basically a write can happen
   -- in any axi state.  AXI has precedence in that catapult write is processed
   -- first at each cycle
  axiWrite: process(ACLK, int_ARESETn)
    -- pragma translate_off
    variable buf : line;
    -- pragma translate_on
    variable i : integer;
    variable useAddr : std_logic_vector(ADDR_WIDTH-1 downto 0);
    variable useAddr2 : std_logic_vector(ADDR_WIDTH-1 downto 0);
  begin
    if (int_ARESETn = '0') then
      AWREADY_reg <= '1';
      AWID_reg <= (others => '0');
      WREADY_reg <= '1';
      BRESP_reg <= AXI4_xRESP_OKAY;
      BVALID_reg <= '0';
      write_state <= axi4w_idle;
      writeAddr <= 0;
      s_wrdy_reg <= '0';
      -- pragma translate_off
      for i in 0 to depth-1 loop 
        mem(i) <= (others => '0');
      end loop;
      -- pragma translate_on
    elsif rising_edge(ACLK) then
      -- When in idle state, catapult and AXI can both initiate writes.
      -- If to the same address, then AXI wins... in this implementation
      if ((s_we = '1') and (write_state = axi4w_idle) and (s_tdone = '0')) then
        mem(to_integer(unsigned(s_waddr))) <= s_dout;
        --write(buf, string'("Slave CAT1 write:mem[0x"));
        --write(buf,  slv2hex(s_waddr));
        --write(buf, string'("]=0x"));
        --write(buf,  slv2hex(s_dout));
        --write(buf, string'(" at T="));
        --write(buf, now);
        --writeline(output, buf);
      end if;
      if ((write_state = axi4w_idle) and (AWVALID = '1')) then
        s_wrdy_reg <= '0';
        AWREADY_reg <= '0';
        AWID_reg <= AWID;
        useAddr := std_logic_vector(shift_right(unsigned(AWADDR) - unsigned(wbase_addr), addrShift));
        -- $display("AWADDR=%d base_address=%d addrShift=%d useAddr=%d at T=%t",
        -- AWADDR, base_address, addrShift, useAddr, $time);
        if (WVALID = '1') then
          -- allow for address and data to be presented in one cycle
          -- Check for the write to be masked
          if (unsigned(WSTRB) /= 0) then -- a byte at a time.  Watch for cwidth much less than DATA_WIDTH
            if (unsigned(useAddr) < depth) then
              for i in 0 to (DATA_WIDTH/8)-1 loop 
                if (WSTRB(i) = '1') then
                  if ((8*i) < cwidth) then
                    if (8*(i+1) <= cwidth) then
                      mem(to_integer(unsigned(useAddr))) (8*(i+1)-1 downto (8*i)) <= WDATA(8*(i+1)-1 downto (8*i));
                    else
                      mem(to_integer(unsigned(useAddr))) (cwidth-1 downto (8*i)) <= WDATA(cwidth-1 downto (8*i));
                    end if;
                  end if;
                end if;
              end loop;
              
              --write(buf, string'("Slave AXI1 write:mem[0x"));
              --write(buf,  slv2hex(useAddr));
              --write(buf, string'("]=0x"));
              --write(buf,  slv2hex(WDATA));
              --write(buf, string'(" at T="));
              --write(buf, now);
              --writeline(output, buf);
            else
              -- pragma translate_off
              write(buf, string'("Error:  Out-of-range AXI memory write access:0x"));
              write(buf,  slv2hex(AWADDR));
              write(buf, string'(" at T="));
              write(buf, now);
              writeline(output, buf);
              -- pragma translate_on
            end if;
          end if;
        end if;
        writeAddr <= to_integer(unsigned(useAddr));
        if ((WLAST = '1') and (WVALID = '1')) then
          write_state <= axi4w_write_done;
          WREADY_reg <= '0';
          BRESP_reg <= AXI4_xRESP_OKAY;
          BVALID_reg <= '1';
        else
          write_state <= axi4w_write;
        end if;
      elsif (write_state = axi4w_write) then
        if (WVALID = '1') then
          useAddr2 := std_logic_vector(to_unsigned(writeAddr+1, useAddr2'length));
          if (unsigned(WSTRB) /= 0) then
            if (unsigned(useAddr2) < depth) then
              for i in 0 to (DATA_WIDTH/8)-1 loop 
                if (WSTRB(i) = '1') then
                  if ((8*i) < cwidth) then
                    if (8*(i+1) <= cwidth) then
                      mem(to_integer(unsigned(useAddr2))) (8*(i+1)-1 downto (8*i)) <= WDATA(8*(i+1)-1 downto (8*i));
                    else
                      mem(to_integer(unsigned(useAddr2))) (cwidth-1 downto (8*i)) <= WDATA(cwidth-1 downto (8*i));
                    end if;
                  end if;
                end if;
              end loop;
              --write(buf, string'("Slave AXI2 write:mem[0x"));
              --write(buf,  slv2hex(useAddr2));
              --write(buf, string'("]=0x"));
              --write(buf,  slv2hex(WDATA));
              --write(buf, string'(" at T="));
              --write(buf, now);
              --writeline(output, buf);
            else 
              -- pragma translate_off
              write(buf, string'("Error:  Out-of-range AXI memory write access:0x"));
              write(buf,  slv2hex(AWADDR));
              write(buf, string'(" at T="));
              write(buf, now);
              writeline(output, buf);
              -- pragma translate_on
            end if;
          end if;
          writeAddr <= to_integer(unsigned(useAddr2));
          if (WLAST = '1') then
            write_state <= axi4w_write_done;
            WREADY_reg <= '0';
            BRESP_reg <= AXI4_xRESP_OKAY;
            BVALID_reg <= '1';
          end if;
        end if;
      elsif (write_state = axi4w_write_done) then
        if (BREADY = '1') then
          AWREADY_reg <= '1';
          WREADY_reg <= '1';
          BRESP_reg <= AXI4_xRESP_OKAY;
          BVALID_reg <= '0';
          write_state <= axi4w_idle;
          s_wrdy_reg <= '1';
        end if;
      else
        s_wrdy_reg <= '1';
      end if;
    end if;
  end process; -- axiWrite

  rCatOutOfOrder <= '1' when (s_re = '1') and
                             (s_rrdy_reg = '1') and
                             (catIsReading = '1') and
                             (next_raddr /= to_integer(unsigned(extCatAddr(s_raddr)))+1)
                  else '0';
  
  -- Catapult read processing
  catRead : process(ACLK, int_ARESETn)
    -- pragma translate_off
    variable buf : line;
    -- pragma translate_on
  begin
    if (int_ARESETn = '0') then
      s_din_reg <= (others => '0');
      s_rrdy_reg <= '0';
      catIsReading <= '0';
      next_raddr <= 0;
    elsif rising_edge(ACLK) then
      -- Catapult has read access to memory
      if (tr_write_done = '1') then
        if ( s_re = '1') then
          --$display("Slave CAT read.  Addr=%x Data=%d T=%t", s_raddr, mem[s_raddr], $time);
          --write(buf, string'("Slave CAT read.  Addr=0x"));
          --write(buf,  slv2hex(s_raddr));
          --write(buf, string'(" Data=0x"));
          --write(buf,  slv2hex(mem(to_integer(unsigned(s_raddr)))));
          --write(buf, string'(" T="));
          --write(buf, now);
          --writeline(output, buf);
          if ((catIsReading = '1') and (rCatOutOfOrder /= '1')) then
            -- Make sure next_addr hasnt incremented off the end
            if (next_raddr < depth) then 
              s_din_reg <= mem(next_raddr);
              next_raddr <= next_raddr+1;
            else
              s_rrdy_reg <= '0';
              catIsReading <= '0';
              next_raddr <= 0;                  
            end if;
          else
            s_din_reg <= mem(to_integer(unsigned(s_raddr)));
            s_rrdy_reg <= '1';
            next_raddr <= to_integer(unsigned(extCatAddr(s_raddr)))+1;
            if ((catIsReading = '1') and (rCatOutOfOrder = '1')) then
              catIsReading <= '0';
            else
              catIsReading <= '1';
            end if;
          end if;
        else
          s_rrdy_reg <= '0';
          catIsReading <= '0';
          next_raddr <= 0;
        end if;
      else
        s_rrdy_reg <= '0';
        catIsReading <= '0';
        next_raddr <= 0;
      end if;
    end if;
  end process;    -- catRead 
  
END rtl;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/ccs_in_v1.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;

PACKAGE ccs_in_pkg_v1 IS

COMPONENT ccs_in_v1
  GENERIC (
    rscid    : INTEGER;
    width    : INTEGER
  );
  PORT (
    idat   : OUT std_logic_vector(width-1 DOWNTO 0);
    dat    : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

END ccs_in_pkg_v1;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY ccs_in_v1 IS
  GENERIC (
    rscid : INTEGER;
    width : INTEGER
  );
  PORT (
    idat  : OUT std_logic_vector(width-1 DOWNTO 0);
    dat   : IN  std_logic_vector(width-1 DOWNTO 0)
  );
END ccs_in_v1;

ARCHITECTURE beh OF ccs_in_v1 IS
BEGIN

  idat <= dat;

END beh;


--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/src/funcs.vhd 

-- a package of attributes that give verification tools a hint about
-- the function being implemented
PACKAGE attributes IS
  ATTRIBUTE CALYPTO_FUNC : string;
  ATTRIBUTE CALYPTO_DATA_ORDER : string;
end attributes;

-----------------------------------------------------------------------
-- Package that declares synthesizable functions needed for RTL output
-----------------------------------------------------------------------

LIBRARY ieee;

use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

PACKAGE funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC;
   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

   FUNCTION maximum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION minimum(arg1, arg2 : INTEGER) RETURN INTEGER;
   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2 : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;
   
-----------------------------------------------------------------
-- logic functions
-----------------------------------------------------------------

   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION or_v (inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;
   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- mux functions
-----------------------------------------------------------------

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC       ) RETURN STD_LOGIC_VECTOR;
   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- latch functions
-----------------------------------------------------------------
   FUNCTION lat_s(dinput: STD_LOGIC       ; clk: STD_LOGIC; doutput: STD_LOGIC       ) RETURN STD_LOGIC;
   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- tristate functions
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC       ; control: STD_LOGIC) RETURN STD_LOGIC;
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION "<" (l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">="(l, r: SIGNED  ) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC;
   FUNCTION ">" (l, r: SIGNED  ) RETURN STD_LOGIC;

   -- RETURN 2 bits (left => lt, right => eq)
   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED;
 
   FUNCTION fabs(arg1: SIGNED  ) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED;
   FUNCTION "**" (l, r: UNSIGNED) RETURN UNSIGNED;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  ;
   FUNCTION "**" (l, r: SIGNED  ) RETURN SIGNED  ;

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-- *_stdar functions use shift functions from std_logic_arith
-----------------------------------------------------------------

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR;

   -----------------------------------------------------------------
   -- *_stdar functions use shift functions from std_logic_arith
   -----------------------------------------------------------------
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED  ;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC;
   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE;
   --FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR;
   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR ;

   FUNCTION ceil_log2(size : NATURAL) return NATURAL;
   FUNCTION bits(size : NATURAL) return NATURAL;    

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR);
   
END funcs;


--------------------------- B O D Y ----------------------------


PACKAGE BODY funcs IS

-----------------------------------------------------------------
-- utility functions
-----------------------------------------------------------------

   FUNCTION TO_STDLOGIC(arg1: BOOLEAN) RETURN STD_LOGIC IS
     BEGIN IF arg1 THEN RETURN '1'; ELSE RETURN '0'; END IF; END;
--   FUNCTION TO_STDLOGIC(arg1: STD_ULOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
--     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: STD_LOGIC_VECTOR(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;
   FUNCTION TO_STDLOGIC(arg1: SIGNED(0 DOWNTO 0)) RETURN STD_LOGIC IS
     BEGIN RETURN arg1(0); END;

   FUNCTION TO_STDLOGICVECTOR(arg1: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
     VARIABLE result: STD_LOGIC_VECTOR(0 DOWNTO 0);
   BEGIN
     result := (0 => arg1);
     RETURN result;
   END;

   FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 > arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION minimum (arg1,arg2: INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 < arg2) THEN
       RETURN(arg1) ;
     ELSE
       RETURN(arg2) ;
     END IF;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;

   FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := input1'LENGTH;
     ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
     ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     --synopsys translate_off
     FOR i IN len-1 DOWNTO 0 LOOP
       result(i) := resolved(input1a(i) & input2a(i));
     END LOOP;
     --synopsys translate_on
     RETURN result;
   END;

   FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED) RETURN UNSIGNED IS
   BEGIN RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

   FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED) RETURN SIGNED IS
   BEGIN RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1), STD_LOGIC_VECTOR(input2))); END;

-----------------------------------------------------------------
-- Logic Functions
-----------------------------------------------------------------

   FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;
   FUNCTION and_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(and_v(inputs, 1)); END;
   FUNCTION or_s (inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(or_v(inputs, 1)); END;
   FUNCTION xor_s(inputs: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
     BEGIN RETURN TO_STDLOGIC(xor_v(inputs, 1)); END;

   FUNCTION and_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result AND inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

   FUNCTION or_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     -- this if is added as a quick fix for a bug in catapult evaluating the loop even if inputs'LENGTH==1
     -- see dts0100971279
     IF icnt2 > 1 THEN
       FOR i IN icnt2-1 DOWNTO 1 LOOP
         inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
         result := result OR inputsx(olenM1 DOWNTO 0);
       END LOOP;
     END IF;
     RETURN result;
   END;

   FUNCTION xor_v(inputs: STD_LOGIC_VECTOR; olen: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT ilen: POSITIVE := inputs'LENGTH;
     CONSTANT ilenM1: POSITIVE := ilen-1; --2.1.6.3
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT ilenMolenM1: INTEGER := ilen-olen-1; --2.1.6.3
     VARIABLE inputsx: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0);
     CONSTANT icnt2: POSITIVE:= inputs'LENGTH/olen;
     VARIABLE result: STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT ilen REM olen = 0 SEVERITY FAILURE;
     --synopsys translate_on
     inputsx := inputs;
     result := inputsx(olenM1 DOWNTO 0);
     FOR i IN icnt2-1 DOWNTO 1 LOOP
       inputsx(ilenMolenM1 DOWNTO 0) := inputsx(ilenM1 DOWNTO olen);
       result := result XOR inputsx(olenM1 DOWNTO 0);
     END LOOP;
     RETURN result;
   END;

-----------------------------------------------------------------
-- Muxes
-----------------------------------------------------------------
   
   FUNCTION mux_sel2_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(1 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 4;
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector( size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "01" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "10" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "11" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel3_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(2 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 8;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000" =>
       result := inputs0(1*size-1 DOWNTO 0*size);
     WHEN "001" =>
       result := inputs0(2*size-1 DOWNTO 1*size);
     WHEN "010" =>
       result := inputs0(3*size-1 DOWNTO 2*size);
     WHEN "011" =>
       result := inputs0(4*size-1 DOWNTO 3*size);
     WHEN "100" =>
       result := inputs0(5*size-1 DOWNTO 4*size);
     WHEN "101" =>
       result := inputs0(6*size-1 DOWNTO 5*size);
     WHEN "110" =>
       result := inputs0(7*size-1 DOWNTO 6*size);
     WHEN "111" =>
       result := inputs0(8*size-1 DOWNTO 7*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel4_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(3 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 16;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "0000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "0001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "0010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "0011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "0100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "0101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "0110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "0111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "1000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "1001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "1010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "1011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "1100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "1101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "1110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "1111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel5_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(4 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 32;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0 );
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "00000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "00001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "00010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "00011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "00100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "00101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "00110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "00111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "01000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "01001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "01010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "01011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "01100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "01101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "01110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "01111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "10000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "10001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "10010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "10011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "10100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "10101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "10110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "10111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "11000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "11001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "11010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "11011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "11100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "11101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "11110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "11111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;
   
   FUNCTION mux_sel6_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR(5 DOWNTO 0))
   RETURN STD_LOGIC_VECTOR IS
     CONSTANT size   : POSITIVE := inputs'LENGTH / 64;
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     VARIABLE result : STD_LOGIC_Vector(size-1 DOWNTO 0);
   BEGIN
     -- for synthesis only
     -- simulation inconsistent with control values 'UXZHLWD'
     CASE sel IS
     WHEN "000000" =>
       result := inputs0( 1*size-1 DOWNTO 0*size);
     WHEN "000001" =>
       result := inputs0( 2*size-1 DOWNTO 1*size);
     WHEN "000010" =>
       result := inputs0( 3*size-1 DOWNTO 2*size);
     WHEN "000011" =>
       result := inputs0( 4*size-1 DOWNTO 3*size);
     WHEN "000100" =>
       result := inputs0( 5*size-1 DOWNTO 4*size);
     WHEN "000101" =>
       result := inputs0( 6*size-1 DOWNTO 5*size);
     WHEN "000110" =>
       result := inputs0( 7*size-1 DOWNTO 6*size);
     WHEN "000111" =>
       result := inputs0( 8*size-1 DOWNTO 7*size);
     WHEN "001000" =>
       result := inputs0( 9*size-1 DOWNTO 8*size);
     WHEN "001001" =>
       result := inputs0( 10*size-1 DOWNTO 9*size);
     WHEN "001010" =>
       result := inputs0( 11*size-1 DOWNTO 10*size);
     WHEN "001011" =>
       result := inputs0( 12*size-1 DOWNTO 11*size);
     WHEN "001100" =>
       result := inputs0( 13*size-1 DOWNTO 12*size);
     WHEN "001101" =>
       result := inputs0( 14*size-1 DOWNTO 13*size);
     WHEN "001110" =>
       result := inputs0( 15*size-1 DOWNTO 14*size);
     WHEN "001111" =>
       result := inputs0( 16*size-1 DOWNTO 15*size);
     WHEN "010000" =>
       result := inputs0( 17*size-1 DOWNTO 16*size);
     WHEN "010001" =>
       result := inputs0( 18*size-1 DOWNTO 17*size);
     WHEN "010010" =>
       result := inputs0( 19*size-1 DOWNTO 18*size);
     WHEN "010011" =>
       result := inputs0( 20*size-1 DOWNTO 19*size);
     WHEN "010100" =>
       result := inputs0( 21*size-1 DOWNTO 20*size);
     WHEN "010101" =>
       result := inputs0( 22*size-1 DOWNTO 21*size);
     WHEN "010110" =>
       result := inputs0( 23*size-1 DOWNTO 22*size);
     WHEN "010111" =>
       result := inputs0( 24*size-1 DOWNTO 23*size);
     WHEN "011000" =>
       result := inputs0( 25*size-1 DOWNTO 24*size);
     WHEN "011001" =>
       result := inputs0( 26*size-1 DOWNTO 25*size);
     WHEN "011010" =>
       result := inputs0( 27*size-1 DOWNTO 26*size);
     WHEN "011011" =>
       result := inputs0( 28*size-1 DOWNTO 27*size);
     WHEN "011100" =>
       result := inputs0( 29*size-1 DOWNTO 28*size);
     WHEN "011101" =>
       result := inputs0( 30*size-1 DOWNTO 29*size);
     WHEN "011110" =>
       result := inputs0( 31*size-1 DOWNTO 30*size);
     WHEN "011111" =>
       result := inputs0( 32*size-1 DOWNTO 31*size);
     WHEN "100000" =>
       result := inputs0( 33*size-1 DOWNTO 32*size);
     WHEN "100001" =>
       result := inputs0( 34*size-1 DOWNTO 33*size);
     WHEN "100010" =>
       result := inputs0( 35*size-1 DOWNTO 34*size);
     WHEN "100011" =>
       result := inputs0( 36*size-1 DOWNTO 35*size);
     WHEN "100100" =>
       result := inputs0( 37*size-1 DOWNTO 36*size);
     WHEN "100101" =>
       result := inputs0( 38*size-1 DOWNTO 37*size);
     WHEN "100110" =>
       result := inputs0( 39*size-1 DOWNTO 38*size);
     WHEN "100111" =>
       result := inputs0( 40*size-1 DOWNTO 39*size);
     WHEN "101000" =>
       result := inputs0( 41*size-1 DOWNTO 40*size);
     WHEN "101001" =>
       result := inputs0( 42*size-1 DOWNTO 41*size);
     WHEN "101010" =>
       result := inputs0( 43*size-1 DOWNTO 42*size);
     WHEN "101011" =>
       result := inputs0( 44*size-1 DOWNTO 43*size);
     WHEN "101100" =>
       result := inputs0( 45*size-1 DOWNTO 44*size);
     WHEN "101101" =>
       result := inputs0( 46*size-1 DOWNTO 45*size);
     WHEN "101110" =>
       result := inputs0( 47*size-1 DOWNTO 46*size);
     WHEN "101111" =>
       result := inputs0( 48*size-1 DOWNTO 47*size);
     WHEN "110000" =>
       result := inputs0( 49*size-1 DOWNTO 48*size);
     WHEN "110001" =>
       result := inputs0( 50*size-1 DOWNTO 49*size);
     WHEN "110010" =>
       result := inputs0( 51*size-1 DOWNTO 50*size);
     WHEN "110011" =>
       result := inputs0( 52*size-1 DOWNTO 51*size);
     WHEN "110100" =>
       result := inputs0( 53*size-1 DOWNTO 52*size);
     WHEN "110101" =>
       result := inputs0( 54*size-1 DOWNTO 53*size);
     WHEN "110110" =>
       result := inputs0( 55*size-1 DOWNTO 54*size);
     WHEN "110111" =>
       result := inputs0( 56*size-1 DOWNTO 55*size);
     WHEN "111000" =>
       result := inputs0( 57*size-1 DOWNTO 56*size);
     WHEN "111001" =>
       result := inputs0( 58*size-1 DOWNTO 57*size);
     WHEN "111010" =>
       result := inputs0( 59*size-1 DOWNTO 58*size);
     WHEN "111011" =>
       result := inputs0( 60*size-1 DOWNTO 59*size);
     WHEN "111100" =>
       result := inputs0( 61*size-1 DOWNTO 60*size);
     WHEN "111101" =>
       result := inputs0( 62*size-1 DOWNTO 61*size);
     WHEN "111110" =>
       result := inputs0( 63*size-1 DOWNTO 62*size);
     WHEN "111111" =>
       result := inputs0( 64*size-1 DOWNTO 63*size);
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_s(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN RETURN TO_STDLOGIC(mux_v(inputs, sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS  --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR(inputs'LENGTH-1 DOWNTO 0) IS inputs;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2 SEVERITY FAILURE;
     --synopsys translate_on
       CASE sel IS
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0( size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1  DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0(size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
       RETURN result;
   END;
--   BEGIN RETURN mux_v(inputs, TO_STDLOGICVECTOR(sel)); END;

   FUNCTION mux_v(inputs: STD_LOGIC_VECTOR; sel : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS --pragma hls_map_to_operator mux
     ALIAS    inputs0: STD_LOGIC_VECTOR( inputs'LENGTH-1 DOWNTO 0) IS inputs;
     ALIAS    sel0   : STD_LOGIC_VECTOR( sel'LENGTH-1 DOWNTO 0 ) IS sel;

     VARIABLE sellen : INTEGER RANGE 2-sel'LENGTH TO sel'LENGTH;
     CONSTANT size   : POSITIVE := inputs'LENGTH / 2;
     CONSTANT olen   : POSITIVE := inputs'LENGTH / 2**sel'LENGTH;
     VARIABLE result : STD_LOGIC_VECTOR(olen-1 DOWNTO 0);
     TYPE inputs_array_type is array(natural range <>) of std_logic_vector( olen - 1 DOWNTO 0);
     VARIABLE inputs_array : inputs_array_type( 2**sel'LENGTH - 1 DOWNTO 0);
   BEGIN
     sellen := sel'LENGTH;
     --synopsys translate_off
     ASSERT inputs'LENGTH = olen * 2**sellen SEVERITY FAILURE;
     sellen := 2-sellen;
     --synopsys translate_on
     CASE sellen IS
     WHEN 1 =>
       CASE sel0(0) IS

       WHEN '1' 
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
            =>
         result := inputs0(  size-1 DOWNTO 0);
       WHEN '0' 
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
            =>
         result := inputs0(2*size-1 DOWNTO size);
       WHEN others =>
         --synopsys translate_off
         result := resolve_std_logic_vector(inputs0( size-1 DOWNTO 0), inputs0( 2*size-1 DOWNTO size));
         --synopsys translate_on
       END CASE;
     WHEN 2 =>
       result := mux_sel2_v(inputs, not sel);
     WHEN 3 =>
       result := mux_sel3_v(inputs, not sel);
     WHEN 4 =>
       result := mux_sel4_v(inputs, not sel);
     WHEN 5 =>
       result := mux_sel5_v(inputs, not sel);
     WHEN 6 =>
       result := mux_sel6_v(inputs, not sel);
     WHEN others =>
       -- synopsys translate_off
       IF(Is_X(sel0)) THEN
         result := (others => 'X');
       ELSE
       -- synopsys translate_on
         FOR i in 0 to 2**sel'LENGTH - 1 LOOP
           inputs_array(i) := inputs0( ((i + 1) * olen) - 1  DOWNTO i*olen);
         END LOOP;
         result := inputs_array(CONV_INTEGER( (UNSIGNED(NOT sel0)) ));
       -- synopsys translate_off
       END IF;
       -- synopsys translate_on
     END CASE;
     RETURN result;
   END;

 
-----------------------------------------------------------------
-- Latches
-----------------------------------------------------------------

   FUNCTION lat_s(dinput: STD_LOGIC; clk: STD_LOGIC; doutput: STD_LOGIC) RETURN STD_LOGIC IS
   BEGIN RETURN mux_s(STD_LOGIC_VECTOR'(doutput & dinput), clk); END;

   FUNCTION lat_v(dinput: STD_LOGIC_VECTOR ; clk: STD_LOGIC; doutput: STD_LOGIC_VECTOR ) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     --synopsys translate_off
     ASSERT dinput'LENGTH = doutput'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN mux_v(doutput & dinput, clk);
   END;

-----------------------------------------------------------------
-- Tri-States
-----------------------------------------------------------------
--   FUNCTION tri_s(dinput: STD_LOGIC; control: STD_LOGIC) RETURN STD_LOGIC IS
--   BEGIN RETURN TO_STDLOGIC(tri_v(TO_STDLOGICVECTOR(dinput), control)); END;
--
--   FUNCTION tri_v(dinput: STD_LOGIC_VECTOR ; control: STD_LOGIC) RETURN STD_LOGIC_VECTOR IS
--     VARIABLE result: STD_LOGIC_VECTOR(dinput'range);
--   BEGIN
--     CASE control IS
--     WHEN '0' | 'L' =>
--       result := (others => 'Z');
--     WHEN '1' | 'H' =>
--       FOR i IN dinput'range LOOP
--         result(i) := to_UX01(dinput(i));
--       END LOOP;
--     WHEN others =>
--       -- synopsys translate_off
--       result := (others => 'X');
--       -- synopsys translate_on
--     END CASE;
--     RETURN result;
--   END;

-----------------------------------------------------------------
-- compare functions returning STD_LOGIC
-- in contrast to the functions returning boolean
-----------------------------------------------------------------

   FUNCTION "=" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;
   FUNCTION "/="(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN or_s(STD_LOGIC_VECTOR(l) xor STD_LOGIC_VECTOR(r)); END;

   FUNCTION "<" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     VARIABLE diff: UNSIGNED(l'LENGTH DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     diff := ('0'&l) - ('0'&r);
     RETURN diff(l'LENGTH);
   END;
   FUNCTION "<"(l, r: SIGNED  ) RETURN STD_LOGIC IS
   BEGIN
     RETURN (UNSIGNED(l) < UNSIGNED(r)) xor (l(l'LEFT) xor r(r'LEFT));
   END;

   FUNCTION "<="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION "<=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(r < l); END;
   FUNCTION ">" (l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">"(l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN r < l; END;
   FUNCTION ">="(l, r: UNSIGNED) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;
   FUNCTION ">=" (l, r: SIGNED  ) RETURN STD_LOGIC IS
     BEGIN RETURN not STD_LOGIC'(l < r); END;

   FUNCTION cmp (l, r: STD_LOGIC_VECTOR) RETURN STD_LOGIC IS
   BEGIN
     --synopsys translate_off
     ASSERT l'LENGTH = r'LENGTH SEVERITY FAILURE;
     --synopsys translate_on
     RETURN not or_s(l xor r);
   END;

-----------------------------------------------------------------
-- Vectorized Overloaded Arithmetic Operators
-----------------------------------------------------------------

   --some functions to placate spyglass
   FUNCTION mult_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a*b;
   END mult_natural;

   FUNCTION div_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a/b;
   END div_natural;

   FUNCTION mod_natural(a,b : NATURAL) RETURN NATURAL IS
   BEGIN
     return a mod b;
   END mod_natural;

   FUNCTION add_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a+b;
   END add_unsigned;

   FUNCTION sub_unsigned(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a-b;
   END sub_unsigned;

   FUNCTION sub_int(a,b : INTEGER) RETURN INTEGER IS
   BEGIN
     return a-b;
   END sub_int;

   FUNCTION concat_0(b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return '0' & b;
   END concat_0;

   FUNCTION concat_uns(a,b : UNSIGNED) RETURN UNSIGNED IS
   BEGIN
     return a&b;
   END concat_uns;

   FUNCTION concat_vect(a,b : STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   BEGIN
     return a&b;
   END concat_vect;





   FUNCTION faccu(arg: UNSIGNED; width: NATURAL) RETURN UNSIGNED IS
     CONSTANT ninps : NATURAL := arg'LENGTH / width;
     ALIAS    arg0  : UNSIGNED(arg'LENGTH-1 DOWNTO 0) IS arg;
     VARIABLE result: UNSIGNED(width-1 DOWNTO 0);
     VARIABLE from  : INTEGER;
     VARIABLE dto   : INTEGER;
   BEGIN
     --synopsys translate_off
     ASSERT arg'LENGTH = width * ninps SEVERITY FAILURE;
     --synopsys translate_on
     result := (OTHERS => '0');
     FOR i IN ninps-1 DOWNTO 0 LOOP
       --result := result + arg0((i+1)*width-1 DOWNTO i*width);
       from := mult_natural((i+1), width)-1; --2.1.6.3
       dto  := mult_natural(i,width); --2.1.6.3
       result := add_unsigned(result , arg0(from DOWNTO dto) );
     END LOOP;
     RETURN result;
   END faccu;

   FUNCTION  fabs (arg1: SIGNED) RETURN UNSIGNED IS
   BEGIN
     CASE arg1(arg1'LEFT) IS
     WHEN '1'
     --synopsys translate_off
          | 'H'
     --synopsys translate_on
       =>
       RETURN UNSIGNED'("0") - UNSIGNED(arg1);
     WHEN '0'
     --synopsys translate_off
          | 'L'
     --synopsys translate_on
       =>
       RETURN UNSIGNED(arg1);
     WHEN others =>
       RETURN resolve_unsigned(UNSIGNED(arg1), UNSIGNED'("0") - UNSIGNED(arg1));
     END CASE;
   END;

   PROCEDURE divmod(l, r: UNSIGNED; rdiv, rmod: OUT UNSIGNED) IS
     CONSTANT llen: INTEGER := l'LENGTH;
     CONSTANT rlen: INTEGER := r'LENGTH;
     CONSTANT llen_plus_rlen: INTEGER := llen + rlen;
     VARIABLE lbuf: UNSIGNED(llen+rlen-1 DOWNTO 0);
     VARIABLE diff: UNSIGNED(rlen DOWNTO 0);
   BEGIN
     --synopsys translate_off
     ASSERT rdiv'LENGTH = llen AND rmod'LENGTH = rlen SEVERITY FAILURE;
     --synopsys translate_on
     lbuf := (others => '0');
     lbuf(llen-1 DOWNTO 0) := l;
     FOR i IN rdiv'range LOOP
       diff := sub_unsigned(lbuf(llen_plus_rlen-1 DOWNTO llen-1) ,(concat_0(r)));
       rdiv(i) := not diff(rlen);
       IF diff(rlen) = '0' THEN
         lbuf(llen_plus_rlen-1 DOWNTO llen-1) := diff;
       END IF;
       lbuf(llen_plus_rlen-1 DOWNTO 1) := lbuf(llen_plus_rlen-2 DOWNTO 0);
     END LOOP;
     rmod := lbuf(llen_plus_rlen-1 DOWNTO llen);
   END divmod;

   FUNCTION "/"  (l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rdiv;
   END "/";

   FUNCTION "MOD"(l, r: UNSIGNED) RETURN UNSIGNED IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(l, r, rdiv, rmod);
     RETURN rmod;
   END;

   FUNCTION "REM"(l, r: UNSIGNED) RETURN UNSIGNED IS
     BEGIN RETURN l MOD r; END;

   FUNCTION "/"  (l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rdiv := UNSIGNED'("0") - rdiv;
     END IF;
     RETURN SIGNED(rdiv); -- overflow problem "1000" / "11"
   END "/";

   FUNCTION "MOD"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
     CONSTANT rnul: UNSIGNED(r'LENGTH-1 DOWNTO 0) := (others => '0');
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     IF rmod /= rnul AND to_X01(l(l'LEFT)) /= to_X01(r(r'LEFT)) THEN
       rmod := UNSIGNED(r) + rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "MOD";

   FUNCTION "REM"(l, r: SIGNED  ) RETURN SIGNED  IS
     VARIABLE rdiv: UNSIGNED(l'LENGTH-1 DOWNTO 0);
     VARIABLE rmod: UNSIGNED(r'LENGTH-1 DOWNTO 0);
   BEGIN
     divmod(fabs(l), fabs(r), rdiv, rmod);
     IF to_X01(l(l'LEFT)) = '1' THEN
       rmod := UNSIGNED'("0") - rmod;
     END IF;
     RETURN SIGNED(rmod);
   END "REM";

   FUNCTION mult_unsigned(l,r : UNSIGNED) return UNSIGNED is
   BEGIN
     return l*r; 
   END mult_unsigned;

   FUNCTION "**" (l, r : UNSIGNED) RETURN UNSIGNED IS
     CONSTANT llen  : NATURAL := l'LENGTH;
     VARIABLE result: UNSIGNED(llen-1 DOWNTO 0);
     VARIABLE fak   : UNSIGNED(llen-1 DOWNTO 0);
   BEGIN
     fak := l;
     result := (others => '0'); result(0) := '1';
     FOR i IN r'reverse_range LOOP
       --was:result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(result & (result*fak)), r(i)));
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR( concat_uns(result , mult_unsigned(result,fak) )), r(i)));

       fak := mult_unsigned(fak , fak);
     END LOOP;
     RETURN result;
   END "**";

   FUNCTION "**" (l, r : SIGNED) RETURN SIGNED IS
     CONSTANT rlen  : NATURAL := r'LENGTH;
     ALIAS    r0    : SIGNED(0 TO r'LENGTH-1) IS r;
     VARIABLE result: SIGNED(l'range);
   BEGIN
     CASE r(r'LEFT) IS
     WHEN '0'
   --synopsys translate_off
          | 'L'
   --synopsys translate_on
     =>
       result := SIGNED(UNSIGNED(l) ** UNSIGNED(r0(1 TO r'LENGTH-1)));
     WHEN '1'
   --synopsys translate_off
          | 'H'
   --synopsys translate_on
     =>
       result := (others => '0');
     WHEN others =>
       result := (others => 'X');
     END CASE;
     RETURN result;
   END "**";

-----------------------------------------------------------------
--               S H I F T   F U C T I O N S
-- negative shift shifts the opposite direction
-----------------------------------------------------------------

   FUNCTION add_nat(arg1 : NATURAL; arg2 : NATURAL ) RETURN NATURAL IS
   BEGIN
     return (arg1 + arg2);
   END;
   
--   FUNCTION UNSIGNED_2_BIT_VECTOR(arg1 : NATURAL; arg2 : NATURAL ) RETURN BIT_VECTOR IS
--   BEGIN
--     return (arg1 + arg2);
--   END;
   
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shl(SIGNED(result), arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
     CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: SIGNED(len-1 DOWNTO 0);
   BEGIN
     result := (others => sbit);
     result(ilenub DOWNTO 0) := arg1;
     result := shr(result, arg2);
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
     --synopsys translate_off
            | 'L'
     --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
     --synopsys translate_off
            | 'H'
     --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
        =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
        =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: SIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl_stdar(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_signed(
           fshr_stdar(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl_stdar(arg1 & '0', '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl_stdar(arg1, arg2, '0', olen); END;
   FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr_stdar(arg1, arg2, '0', olen); END;

   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;
   FUNCTION fshr_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN fshr_stdar(arg1, arg2, arg1(arg1'LEFT), olen); END;


   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     --SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: NATURAL range 1 TO len;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => '0');
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         --was:temp(i2+sw) := result(i2);
         temp_idx := add_nat(i2,sw);
         temp(temp_idx) := result(i2);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT ilen: INTEGER := arg1'LENGTH;
     CONSTANT olenM1: INTEGER := olen-1; --2.1.6.3
     CONSTANT len: INTEGER := maximum(ilen, olen);
     VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
     VARIABLE temp: UNSIGNED(len-1 DOWNTO 0);
     SUBTYPE  sw_range IS NATURAL range 1 TO len;
     VARIABLE sw: sw_range;
     VARIABLE result_idx : INTEGER; --2.1.6.3
   BEGIN
     sw := 1;
     result := (others => sbit);
     result(ilen-1 DOWNTO 0) := arg1;
     FOR i IN arg2'reverse_range LOOP
       temp := (others => sbit);
       FOR i2 IN len-1-sw DOWNTO 0 LOOP
         -- was: temp(i2) := result(i2+sw);
         result_idx := add_nat(i2,sw);
         temp(i2) := result(result_idx);
       END LOOP;
       result := UNSIGNED(mux_v(STD_LOGIC_VECTOR(concat_uns(result,temp)), arg2(i)));
       sw := minimum(mult_natural(sw,2), len);
     END LOOP;
     RETURN result(olenM1 DOWNTO 0);
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
     ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
     CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others=>'0');
     arg1x_pad(arg1l+1) := sbit;
     arg1x_pad(arg1l downto 0) := arg1x;
     IF arg2l = 0 THEN
       RETURN fshr(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
     -- ELSIF arg1l = 0 THEN
     --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshl(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
           fshr(arg1x_pad(arg1l+1 DOWNTO 1), not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
         );
         --synopsys translate_on
         RETURN result;
       END CASE;
     END IF;
   END;

   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
     CONSTANT arg2l: INTEGER := arg2'LENGTH - 1;
     ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
     VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
   BEGIN
     result := (others => '0');
     IF arg2l = 0 THEN
       RETURN fshl(arg1, UNSIGNED(arg2x), olen);
     ELSE
       CASE arg2x(arg2l) IS
       WHEN '0'
       --synopsys translate_off
            | 'L'
       --synopsys translate_on
       =>
         RETURN fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);

       WHEN '1'
       --synopsys translate_off
            | 'H'
       --synopsys translate_on
       =>
         RETURN fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen);
       WHEN others =>
         --synopsys translate_off
         result := resolve_unsigned(
           fshr(arg1, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen),
           fshl(arg1 & '0', not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), olen)
         );
         --synopsys translate_on
	 return result;
       END CASE;
     END IF;
   END;

   FUNCTION fshl(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;
   FUNCTION fshl(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshl(arg1, arg2, '0', olen); END;
   FUNCTION fshr(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE) RETURN UNSIGNED IS
     BEGIN RETURN fshr(arg1, arg2, '0', olen); END;

   FUNCTION fshl(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshl(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshl(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;
   FUNCTION fshr(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE) RETURN SIGNED   IS
     BEGIN RETURN SIGNED(fshr(UNSIGNED(arg1), arg2, arg1(arg1'LEFT), olen)); END;


   FUNCTION frot(arg1: STD_LOGIC_VECTOR; arg2: STD_LOGIC_VECTOR; signd2: BOOLEAN; sdir: INTEGER range -1 TO 1) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len: INTEGER := arg1'LENGTH;
     VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     VARIABLE temp: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     SUBTYPE sw_range IS NATURAL range 0 TO len-1;
     VARIABLE sw: sw_range;
     VARIABLE temp_idx : INTEGER; --2.1.6.3
   BEGIN
     result := (others=>'0');
     result := arg1;
     sw := sdir MOD len;
     FOR i IN arg2'reverse_range LOOP
       EXIT WHEN sw = 0;
       IF signd2 AND i = arg2'LEFT THEN 
         sw := sub_int(len,sw); 
       END IF;
       -- temp := result(len-sw-1 DOWNTO 0) & result(len-1 DOWNTO len-sw)
       FOR i2 IN len-1 DOWNTO 0 LOOP
         --was: temp((i2+sw) MOD len) := result(i2);
         temp_idx := add_nat(i2,sw) MOD len;
         temp(temp_idx) := result(i2);
       END LOOP;
       result := mux_v(STD_LOGIC_VECTOR(concat_vect(result,temp)), arg2(i));
       sw := mod_natural(mult_natural(sw,2), len);
     END LOOP;
     RETURN result;
   END frot;

   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: UNSIGNED) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), FALSE, -1); END;
   FUNCTION frol(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, 1); END;
   FUNCTION fror(arg1: STD_LOGIC_VECTOR; arg2: SIGNED  ) RETURN STD_LOGIC_VECTOR IS
     BEGIN RETURN frot(arg1, STD_LOGIC_VECTOR(arg2), TRUE, -1); END;

-----------------------------------------------------------------
-- indexing functions: LSB always has index 0
-----------------------------------------------------------------

   FUNCTION readindex(vec: STD_LOGIC_VECTOR; index: INTEGER                 ) RETURN STD_LOGIC IS
     CONSTANT len : INTEGER := vec'LENGTH;
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
   BEGIN
     IF index >= len OR index < 0 THEN
       RETURN 'X';
     END IF;
     RETURN vec0(index);
   END;

   FUNCTION readslice(vec: STD_LOGIC_VECTOR; index: INTEGER; width: POSITIVE) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     CONSTANT indexPwidthM1 : INTEGER := index+width-1; --2.1.6.3
     ALIAS    vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS vec;
     CONSTANT xxx : STD_LOGIC_VECTOR(width-1 DOWNTO 0) := (others => 'X');
   BEGIN
     IF index+width > len OR index < 0 THEN
       RETURN xxx;
     END IF;
     RETURN vec0(indexPwidthM1 DOWNTO index);
   END;

   FUNCTION writeindex(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC       ; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
     CONSTANT len : INTEGER := vec'LENGTH;
     VARIABLE vec0: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
     CONSTANT xxx : STD_LOGIC_VECTOR(len-1 DOWNTO 0) := (others => 'X');
   BEGIN
     vec0 := vec;
     IF index >= len OR index < 0 THEN
       RETURN xxx;
     END IF;
     vec0(index) := dinput;
     RETURN vec0;
   END;

   FUNCTION n_bits(p: NATURAL) RETURN POSITIVE IS
     VARIABLE n_b : POSITIVE;
     VARIABLE p_v : NATURAL;
   BEGIN
     p_v := p;
     FOR i IN 1 TO 32 LOOP
       p_v := div_natural(p_v,2);
       n_b := i;
       EXIT WHEN (p_v = 0);
     END LOOP;
     RETURN n_b;
   END;


--   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; index: INTEGER) RETURN STD_LOGIC_VECTOR IS
--
--     CONSTANT vlen: INTEGER := vec'LENGTH;
--     CONSTANT ilen: INTEGER := dinput'LENGTH;
--     CONSTANT max_shift: INTEGER := vlen-ilen;
--     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
--     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
--     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
--     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
--     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
--     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
--   BEGIN
--     inp := (others => '0');
--     mask := (others => '0');
--
--     IF index > max_shift OR index < 0 THEN
--       RETURN xxx;
--     END IF;
--
--     shift := CONV_UNSIGNED(index, shift'LENGTH);
--     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
--     mask(ilen-1 DOWNTO 0) := ones;
--     inp := fshl(inp, shift, vlen);
--     mask := fshl(mask, shift, vlen);
--     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
--     RETURN vec0;
--   END;

   FUNCTION writeslice(vec: STD_LOGIC_VECTOR; dinput: STD_LOGIC_VECTOR; enable: STD_LOGIC_VECTOR; byte_width: INTEGER;  index: INTEGER) RETURN STD_LOGIC_VECTOR IS

     type enable_matrix is array (0 to enable'LENGTH-1 ) of std_logic_vector(byte_width-1 downto 0);
     CONSTANT vlen: INTEGER := vec'LENGTH;
     CONSTANT ilen: INTEGER := dinput'LENGTH;
     CONSTANT max_shift: INTEGER := vlen-ilen;
     CONSTANT ones: UNSIGNED(ilen-1 DOWNTO 0) := (others => '1');
     CONSTANT xxx : STD_LOGIC_VECTOR(vlen-1 DOWNTO 0) := (others => 'X');
     VARIABLE shift : UNSIGNED(n_bits(max_shift)-1 DOWNTO 0);
     VARIABLE vec0: STD_LOGIC_VECTOR(vlen-1 DOWNTO 0);
     VARIABLE inp: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE mask2: UNSIGNED(vlen-1 DOWNTO 0);
     VARIABLE enables: enable_matrix;
     VARIABLE cat_enables: STD_LOGIC_VECTOR(ilen-1 DOWNTO 0 );
     VARIABLE lsbi : INTEGER;
     VARIABLE msbi : INTEGER;

   BEGIN
     cat_enables := (others => '0');
     lsbi := 0;
     msbi := byte_width-1;
     inp := (others => '0');
     mask := (others => '0');

     IF index > max_shift OR index < 0 THEN
       RETURN xxx;
     END IF;

     --initialize enables
     for i in 0 TO (enable'LENGTH-1) loop
       enables(i)  := (others => enable(i));
       cat_enables(msbi downto lsbi) := enables(i) ;
       lsbi := msbi+1;
       msbi := msbi+byte_width;
     end loop;


     shift := CONV_UNSIGNED(index, shift'LENGTH);
     inp(ilen-1 DOWNTO 0) := UNSIGNED(dinput);
     mask(ilen-1 DOWNTO 0) := UNSIGNED((STD_LOGIC_VECTOR(ones) AND cat_enables));
     inp := fshl(inp, shift, vlen);
     mask := fshl(mask, shift, vlen);
     vec0 := (vec and (not STD_LOGIC_VECTOR(mask))) or STD_LOGIC_VECTOR(inp);
     RETURN vec0;
   END;


   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;
   
   FUNCTION bits(size : NATURAL) return NATURAL is
   begin
     return ceil_log2(size);
   END;

   PROCEDURE csa(a, b, c: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH) xor conv_std_logic_vector(c, s'LENGTH);
     cout := ( (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH)) or (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) or (conv_std_logic_vector(b, cout'LENGTH) and conv_std_logic_vector(c, cout'LENGTH)) );
   END PROCEDURE csa;

   PROCEDURE csha(a, b: IN INTEGER; s, cout: OUT STD_LOGIC_VECTOR) IS
   BEGIN
     s    := conv_std_logic_vector(a, s'LENGTH) xor conv_std_logic_vector(b, s'LENGTH);
     cout := (conv_std_logic_vector(a, cout'LENGTH) and conv_std_logic_vector(b, cout'LENGTH));
   END PROCEDURE csha;

END funcs;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_comps.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_comps IS
 
FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER;
FUNCTION ceil_log2(size : NATURAL) return NATURAL;
 

COMPONENT mgc_not
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_and
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nand
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_or
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_nor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_xnor
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux
  GENERIC (
    width  :  NATURAL;
    ctrlw  :  NATURAL;
    p2ctrlw : NATURAL := 0
  );
  PORT (
    a: in  std_logic_vector(width*(2**ctrlw) - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw            - 1 DOWNTO 0);
    z: out std_logic_vector(width            - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mux1hot
  GENERIC (
    width  : NATURAL;
    ctrlw  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ctrlw - 1 DOWNTO 0);
    c: in  std_logic_vector(ctrlw       - 1 DOWNTO 0);
    z: out std_logic_vector(width       - 1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_reg_pos
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;  -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL  -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_reg_neg
  GENERIC (
    width  : NATURAL;
    has_a_rst : NATURAL;  -- 0 to 1
    a_rst_on  : NATURAL;  -- 0 to 1
    has_s_rst : NATURAL;  -- 0 to 1
    s_rst_on  : NATURAL;   -- 0 to 1
    has_enable : NATURAL; -- 0 to 1
    enable_on  : NATURAL -- 0 to 1
  );
  PORT (
    clk: in  std_logic;
    d  : in  std_logic_vector(width-1 DOWNTO 0);
    z  : out std_logic_vector(width-1 DOWNTO 0);
    sync_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    sync_rst : in std_logic;
    async_rst_val : in std_logic_vector(width-1 DOWNTO 0);
    async_rst : in std_logic;
    en : in std_logic
  );
END COMPONENT;

COMPONENT mgc_generic_reg
  GENERIC(
   width: natural := 8;
   ph_clk: integer range 0 to 1 := 1; -- clock polarity, 1=rising_edge
   ph_en: integer range 0 to 1 := 1;
   ph_a_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   ph_s_rst: integer range 0 to 1 := 1;   --  0 to 1 IGNORED
   a_rst_used: integer range 0 to 1 := 1;
   s_rst_used: integer range 0 to 1 := 0;
   en_used: integer range 0 to 1 := 1
  );
  PORT(
   d: std_logic_vector(width-1 downto 0);
   clk: in std_logic;
   en: in std_logic;
   a_rst: in std_logic;
   s_rst: in std_logic;
   q: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_equal
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a : in  std_logic_vector(width-1 DOWNTO 0);
    b : in  std_logic_vector(width-1 DOWNTO 0);
    eq: out std_logic;
    ne: out std_logic
  );
END COMPONENT;

COMPONENT mgc_shift_l
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rot
  GENERIC (
    width  : NATURAL;
    width_s: NATURAL;
    signd_s: NATURAL;      -- 0:unsigned 1:signed
    sleft  : NATURAL;      -- 0:right 1:left;
    log2w  : NATURAL := 0; -- LOG2(width)
    l2wp2  : NATURAL := 0  --2**LOG2(width)
  );
  PORT (
    a : in  std_logic_vector(width  -1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width  -1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_sub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_ci
  GENERIC (
    width_a : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width_a, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width_a, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width_a,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width_a,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_addc
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add3
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_c : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_c : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    c: in  std_logic_vector(ifeqsel(width_c,0,width,width_c)-1 DOWNTO 0);
    d: in  std_logic_vector(0 DOWNTO 0);
    e: in  std_logic_vector(0 DOWNTO 0);
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_add_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_sub_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addc_pipe
  GENERIC (
     width_a : natural := 16;
     signd_a : integer range 0 to 1 := 0;
     width_b : natural := 3;
     signd_b : integer range 0 to 1 := 0;
     width_z : natural := 18;
     ph_clk : integer range 0 to 1 := 1;
     ph_en : integer range 0 to 1 := 1;
     ph_a_rst : integer range 0 to 1 := 1;
     ph_s_rst : integer range 0 to 1 := 1;
     n_outreg : natural := 2;
     stages : natural := 2; -- Default value is minimum required value
     a_rst_used: integer range 0 to 1 := 1;
     s_rst_used: integer range 0 to 1 := 0;
     en_used: integer range 0 to 1 := 1
     );
  PORT(
     a: in std_logic_vector(width_a-1 downto 0);
     b: in std_logic_vector(width_b-1 downto 0);
     c: in std_logic_vector(0 downto 0);
     clk: in std_logic;
     en: in std_logic;
     a_rst: in std_logic;
     s_rst: in std_logic;
     z: out std_logic_vector(width_z-1 downto 0)
     );
END COMPONENT;

COMPONENT mgc_addsub
  GENERIC (
    width   : NATURAL; 
    signd_a : NATURAL := 0;
    width_b : NATURAL := 0; -- if == 0 use width, compatiability with versions < 2005a
    signd_b : NATURAL := 0;
    width_z : NATURAL := 0  -- if == 0 use width, compatiability with versions < 2005a
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    b: in  std_logic_vector(ifeqsel(width_b,0,width,width_b)-1 DOWNTO 0);
    add: in  std_logic;
    z: out std_logic_vector(ifeqsel(width_z,0,width,width_z)-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_accu
  GENERIC (
    width  : NATURAL;
    ninps  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width*ninps-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_abs
  GENERIC (
    width  : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width-1 DOWNTO 0);
    z: out std_logic_vector(width-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_fast
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_z : NATURAL    -- <= width_a + width_b
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul_pipe
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;   -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2  : NATURAL;
    add_d2  : NATURAL
  );
  PORT (
    a   : in  std_logic_vector(width_a-1 DOWNTO 0);
    b   : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2  : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c   : in  std_logic_vector(width_c-1 DOWNTO 0);
    d   : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2  : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst : in  std_logic_vector(width_e-1 DOWNTO 0);
    z   : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2add1_pipe
  GENERIC (
    gentype : NATURAL;
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_b2 : NATURAL;
    signd_b2 : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_d2 : NATURAL;
    signd_d2 : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c + width_d)+1
    isadd   : NATURAL;
    add_b2   : NATURAL;
    add_d2   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    b2     : in  std_logic_vector(width_b2-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    d2     : in  std_logic_vector(width_d2-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_e-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL
  );
  PORT (
    a:   in  std_logic_vector(width_a-1 DOWNTO 0);
    b:   in  std_logic_vector(width_b-1 DOWNTO 0);
    c:   in  std_logic_vector(width_c-1 DOWNTO 0);
    cst: in  std_logic_vector(width_cst-1 DOWNTO 0);
    d:   in  std_logic_vector(width_d-1 DOWNTO 0);
    z:   out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_muladd1_pipe
  -- operation is z = a * (b + d) + c + cst
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_cst : NATURAL;
    signd_cst : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c, width_cst)+1
    add_axb : NATURAL;
    add_c   : NATURAL;
    add_d   : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    c     : in  std_logic_vector(width_c-1 DOWNTO 0);
    cst   : in  std_logic_vector(width_cst-1 DOWNTO 0);
    d     : in  std_logic_vector(width_d-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mulacc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mul2acc_pipe
  GENERIC (
    width_a : NATURAL;
    signd_a : NATURAL;
    width_b : NATURAL;
    signd_b : NATURAL;
    width_c : NATURAL;
    signd_c : NATURAL;
    width_d : NATURAL;
    signd_d : NATURAL;
    width_e : NATURAL;
    signd_e : NATURAL;
    width_z : NATURAL;    -- <= max(width_a + width_b, width_c)+1
    add_cxd : NATURAL;
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 
  );
  PORT (
    a         : in  std_logic_vector(width_a-1 DOWNTO 0);
    b         : in  std_logic_vector(width_b-1 DOWNTO 0);
    c         : in  std_logic_vector(width_c-1 DOWNTO 0);
    d         : in  std_logic_vector(width_d-1 DOWNTO 0);
    e         : in  std_logic_vector(width_e-1 DOWNTO 0);
    load      : in  std_logic;
    datavalid : in  std_logic;
    clk       : in  std_logic;
    en        : in  std_logic;
    a_rst     : in  std_logic;
    s_rst     : in  std_logic;
    z         : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_div
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_a-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_mod
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_rem
  GENERIC (
    width_a : NATURAL;
    width_b : NATURAL;
    signd   : NATURAL
  );
  PORT (
    a: in  std_logic_vector(width_a-1 DOWNTO 0);
    b: in  std_logic_vector(width_b-1 DOWNTO 0);
    z: out std_logic_vector(width_b-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_csa
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     c: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_csha
  GENERIC (
     width : NATURAL
  );
  PORT (
     a: in std_logic_vector(width-1 downto 0);
     b: in std_logic_vector(width-1 downto 0);
     s: out std_logic_vector(width-1 downto 0);
     cout: out std_logic_vector(width-1 downto 0)
  );
END COMPONENT;

COMPONENT mgc_rom
    GENERIC (
      rom_id : natural := 1;
      size : natural := 33;
      width : natural := 32
      );
    PORT (
      data_in : std_logic_vector((size*width)-1 downto 0);
      addr : std_logic_vector(ceil_log2(size)-1 downto 0);
      data_out : out std_logic_vector(width-1 downto 0)
    );
END COMPONENT;

END mgc_comps;

PACKAGE BODY mgc_comps IS
 
   FUNCTION ceil_log2(size : NATURAL) return NATURAL is
     VARIABLE cnt : NATURAL;
     VARIABLE res : NATURAL;
   begin
     cnt := 1;
     res := 0;
     while (cnt < size) loop
       res := res + 1;
       cnt := 2 * cnt;
     end loop;
     return res;
   END;

   FUNCTION ifeqsel(arg1, arg2, seleq, selne : INTEGER) RETURN INTEGER IS
   BEGIN
     IF(arg1 = arg2) THEN
       RETURN(seleq) ;
     ELSE
       RETURN(selne) ;
     END IF;
   END;
 
END mgc_comps;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/hls_pkgs/mgc_comps_src/mgc_mul_pipe_beh.vhd 

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_mul_pipe IS
  GENERIC (
    width_a       : NATURAL;
    signd_a       : NATURAL;
    width_b       : NATURAL;
    signd_b       : NATURAL;
    width_z       : NATURAL; -- <= width_a + width_b
    clock_edge    : NATURAL; -- 0 to 1
    enable_active : NATURAL; -- 0 to 1
    a_rst_active  : NATURAL; -- 0 to 1 IGNORED
    s_rst_active  : NATURAL; -- 0 to 1 IGNORED
    stages        : NATURAL;    
    n_inreg       : NATURAL := 0 -- default for backwards compatability 

  );
  PORT (
    a     : in  std_logic_vector(width_a-1 DOWNTO 0);
    b     : in  std_logic_vector(width_b-1 DOWNTO 0);
    clk   : in  std_logic;
    en    : in  std_logic;
    a_rst : in  std_logic;
    s_rst : in  std_logic;
    z     : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_mul_pipe;

LIBRARY IEEE;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_mul_pipe IS
  TYPE reg_array_type is array(natural range<>) of std_logic_vector(width_z-1 DOWNTO 0); 
  SIGNAL xz : std_logic_vector(width_a+width_b DOWNTO 0);

--MF Added pipelined input
    signal a_f     : STD_LOGIC_VECTOR(width_a-1 downto 0); 
    signal b_f     : STD_LOGIC_VECTOR(width_b-1 downto 0);
   type a_array is array (natural range <>) of STD_LOGIC_VECTOR(width_a-1 downto 0);
   type b_array is array (natural range <>) of STD_LOGIC_VECTOR(width_b-1 downto 0);
BEGIN
  n_inreg_gt_0: if n_inreg > 0 generate
    GENPOS_INREG: IF clock_edge = 1 GENERATE
     I0: process(clk)
        variable a_in_reg: a_array(n_inreg-1 downto 0);
        variable b_in_reg: b_array(n_inreg-1 downto 0);
      begin
        if (clk'event and clk = '1' ) then
          if (conv_integer(en) = enable_active) then
            for i in n_inreg - 2 downto 0 loop
              a_in_reg(i+1) := a_in_reg(i);
              b_in_reg(i+1) := b_in_reg(i);
            end loop;                                                                                                                             
            a_in_reg(0) := a;
            b_in_reg(0) := b;

            a_f <= a_in_reg(n_inreg-1);             
            b_f <= b_in_reg(n_inreg-1);    
                                                   
          end if;
        end if;
      end process;
    END GENERATE;
  
   GENNEG_INREG: IF clock_edge = 0 GENERATE
     I0: process(clk)
        variable a_in_reg: a_array(n_inreg-1 downto 0);
        variable b_in_reg: b_array(n_inreg-1 downto 0);
      begin
        if (clk'event and clk = '0' ) then
          if (conv_integer(en) = enable_active) then
            for i in n_inreg - 2 downto 0 loop
              a_in_reg(i+1) := a_in_reg(i);
              b_in_reg(i+1) := b_in_reg(i);
            end loop;                                                                                                                             
            a_in_reg(0) := a;
            b_in_reg(0) := b;            
                                 
            a_f <= a_in_reg(n_inreg-1);             
            b_f <= b_in_reg(n_inreg-1);
                                                        
          end if;
        end if;
      end process;
    END GENERATE;
  END GENERATE;

  n_inreg_eq_0: if n_inreg = 0 generate
    a_f <= a;
    b_f <= b;
  end generate n_inreg_eq_0;

  xz <= '0'&(unsigned(a_f) * unsigned(b_f)) WHEN signd_a = 0 AND signd_b = 0 ELSE
            (  signed(a_f) * unsigned(b_f)) WHEN signd_a = 1 AND signd_b = 0 ELSE
            (unsigned(a_f) *   signed(b_f)) WHEN signd_a = 0 AND signd_b = 1 ELSE
        '0'&(  signed(a_f) *   signed(b_f));

  GENPOS: IF clock_edge = 1 GENERATE
    PROCESS (clk)
    VARIABLE reg_array: reg_array_type(stages-2 DOWNTO 0);
    BEGIN
      IF ( clk'EVENT AND clk = '1') THEN
        IF ( conv_integer(en) = enable_active) THEN
          FOR I IN stages-2 DOWNTO 1 LOOP
            reg_array(I) := reg_array(I-1);
          END LOOP;
          reg_array(0) := xz(width_z-1 DOWNTO 0);
          z <= reg_array(stages-2);
        END IF;
      END IF;
    END PROCESS;
  END GENERATE;

  GENNEG: IF clock_edge = 0 GENERATE
    PROCESS (clk)
    VARIABLE reg_array: reg_array_type(stages-2 DOWNTO 0);
    BEGIN
      IF ( clk'EVENT AND clk = '0') THEN
        IF ( conv_integer(en) = enable_active) THEN
          FOR I IN stages-2 DOWNTO 1 LOOP
            reg_array(I) := reg_array(I-1);
          END LOOP;
          reg_array(0) := xz(width_z-1 DOWNTO 0);
          z <= reg_array(stages-2);
        END IF;
      END IF;
    END PROCESS;
  END GENERATE;
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_comps_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;

PACKAGE mgc_shift_comps_v5 IS

COMPONENT mgc_shift_l_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_r_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_bl_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

COMPONENT mgc_shift_br_v5
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END COMPONENT;

END mgc_shift_comps_v5;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_bl_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_bl_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_bl_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_bl_v5 IS

  FUNCTION resolve_std_logic_vector(input1: STD_LOGIC_VECTOR; input2: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
    CONSTANT len: INTEGER := input1'LENGTH;
    ALIAS input1a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input1;
    ALIAS input2a: STD_LOGIC_VECTOR(len-1 DOWNTO 0) IS input2;
    VARIABLE result: STD_LOGIC_VECTOR(len-1 DOWNTO 0);
  BEGIN
    result := (others => '0');
    --synopsys translate_off
    FOR i IN len-1 DOWNTO 0 LOOP
      result(i) := resolved(input1a(i) & input2a(i));
    END LOOP;
    --synopsys translate_on
    RETURN result;
  END;

  FUNCTION resolve_unsigned(input1: UNSIGNED; input2: UNSIGNED)
  RETURN UNSIGNED IS
  BEGIN
    RETURN UNSIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1),
                                             STD_LOGIC_VECTOR(input2)));
  END;

  FUNCTION resolve_signed(input1: SIGNED; input2: SIGNED)
  RETURN SIGNED IS
  BEGIN
    RETURN SIGNED(resolve_std_logic_vector(STD_LOGIC_VECTOR(input1),
                                           STD_LOGIC_VECTOR(input2)));
  END;

  FUNCTION "not"(arg1: UNSIGNED) RETURN UNSIGNED IS
    BEGIN RETURN UNSIGNED(not STD_LOGIC_VECTOR(arg1)); END;

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshr_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shr(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshr_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shr(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

 FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
    ALIAS    arg1x: UNSIGNED(arg1l DOWNTO 0) IS arg1;
    CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
    ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
    VARIABLE arg1x_pad: UNSIGNED(arg1l+1 DOWNTO 0);
    VARIABLE result: UNSIGNED(olen-1 DOWNTO 0);
  BEGIN
    result := (others=>'0');
    arg1x_pad(arg1l+1) := sbit;
    arg1x_pad(arg1l downto 0) := arg1x;
    IF arg2l = 0 THEN
      RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
    -- ELSIF arg1l = 0 THEN
    --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
    ELSE
      CASE arg2x(arg2l) IS
      WHEN '0'
    --synopsys translate_off
           | 'L'
    --synopsys translate_on
      =>
        RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN '1'
    --synopsys translate_off
           | 'H'
    --synopsys translate_on
      =>
        RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN others =>
        --synopsys translate_off
        result := resolve_unsigned(
          fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
          fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
        );
        --synopsys translate_on
        RETURN result;
      END CASE;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: SIGNED  ; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT arg1l: NATURAL := arg1'LENGTH - 1;
    ALIAS    arg1x: SIGNED(arg1l DOWNTO 0) IS arg1;
    CONSTANT arg2l: NATURAL := arg2'LENGTH - 1;
    ALIAS    arg2x: SIGNED(arg2l DOWNTO 0) IS arg2;
    VARIABLE arg1x_pad: SIGNED(arg1l+1 DOWNTO 0);
    VARIABLE result: SIGNED(olen-1 DOWNTO 0);
  BEGIN
    result := (others=>'0');
    arg1x_pad(arg1l+1) := sbit;
    arg1x_pad(arg1l downto 0) := arg1x;
    IF arg2l = 0 THEN
      RETURN fshr_stdar(arg1x_pad, UNSIGNED(arg2x), sbit, olen);
    -- ELSIF arg1l = 0 THEN
    --   RETURN fshl(sbit & arg1x, arg2x, sbit, olen);
    ELSE
      CASE arg2x(arg2l) IS
      WHEN '0'
      --synopsys translate_off
           | 'L'
      --synopsys translate_on
      =>
        RETURN fshl_stdar(arg1x_pad, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN '1'
      --synopsys translate_off
           | 'H'
      --synopsys translate_on
      =>
        RETURN fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen);
      WHEN others =>
        --synopsys translate_off
        result := resolve_signed(
          fshl_stdar(arg1x, UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit,  olen),
          fshr_stdar(arg1x_pad(arg1l+1 DOWNTO 1), '0' & not UNSIGNED(arg2x(arg2l-1 DOWNTO 0)), sbit, olen)
        );
        --synopsys translate_on
        RETURN result;
      END CASE;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: SIGNED  ; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: SIGNED  ; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), signed(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), signed(s), width_z));
  END GENERATE;
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.vhd 
LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY mgc_shift_l_v5 IS
  GENERIC (
    width_a: NATURAL;
    signd_a: NATURAL;
    width_s: NATURAL;
    width_z: NATURAL
  );
  PORT (
    a : in  std_logic_vector(width_a-1 DOWNTO 0);
    s : in  std_logic_vector(width_s-1 DOWNTO 0);
    z : out std_logic_vector(width_z-1 DOWNTO 0)
  );
END mgc_shift_l_v5;

LIBRARY ieee;

USE ieee.std_logic_arith.all;

ARCHITECTURE beh OF mgc_shift_l_v5 IS

  FUNCTION maximum (arg1,arg2: INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1 > arg2) THEN
      RETURN(arg1) ;
    ELSE
      RETURN(arg2) ;
    END IF;
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN UNSIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: UNSIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(result, arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED; arg2: UNSIGNED; sbit: STD_LOGIC; olen: POSITIVE) RETURN SIGNED IS
    CONSTANT ilen: INTEGER := arg1'LENGTH;
    CONSTANT olenM1: INTEGER := olen-1; -- 2.1.6.3
    CONSTANT ilenub: INTEGER := arg1'LENGTH-1;
    CONSTANT len: INTEGER := maximum(ilen, olen);
    VARIABLE result: SIGNED(len-1 DOWNTO 0);
  BEGIN
    result := (others => sbit);
    result(ilenub DOWNTO 0) := arg1;
    result := shl(SIGNED(result), arg2);
    RETURN result(olenM1 DOWNTO 0);
  END;

  FUNCTION fshl_stdar(arg1: UNSIGNED; arg2: UNSIGNED; olen: POSITIVE)
  RETURN UNSIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, '0', olen);
  END;

  FUNCTION fshl_stdar(arg1: SIGNED  ; arg2: UNSIGNED; olen: POSITIVE)
  RETURN SIGNED IS
  BEGIN
    RETURN fshl_stdar(arg1, arg2, arg1(arg1'LEFT), olen);
  END;

BEGIN
UNSGNED:  IF signd_a = 0 GENERATE
    z <= std_logic_vector(fshl_stdar(unsigned(a), unsigned(s), width_z));
  END GENERATE;
SGNED:  IF signd_a /= 0 GENERATE
    z <= std_logic_vector(fshl_stdar(  signed(a), unsigned(s), width_z));
  END GENERATE;
END beh;

--------> /opt/mentorgraphics/Catapult_10.5c/Mgc_home/pkgs/ccs_xilinx/hdl/BLOCK_2R1W_RBW.vhd 
-- Memory Type:            BLOCK
-- Operating Mode:         Unknown Memory Type
-- Clock Mode:             Single Clock
-- 
-- RTL Code RW Resolution: RBW
-- Catapult RW Resolution: RBW
-- 
-- HDL Work Library:       Xilinx_RAMS_lib
-- Component Name:         BLOCK_2R1W_RBW
-- Latency = 1:            RAM with no registers on inputs or outputs
--         = 2:            adds embedded register on RAM output
--         = 3:            adds fabric registers to non-clock input RAM pins
--         = 4:            adds fabric register to output (driven by embedded register from latency=2)

LIBRARY ieee;

  USE ieee.std_logic_1164.all;
  USE ieee.numeric_std.all;
PACKAGE BLOCK_2R1W_RBW_pkg IS
  COMPONENT BLOCK_2R1W_RBW IS
  GENERIC (
    addr_width : integer := 8 ;
    data_width : integer := 7 ;
    depth : integer := 256 ;
    latency : integer := 1 
    
  );
  PORT (
    adra : in std_logic_vector(addr_width-1 downto 0) ;
    adrb : in std_logic_vector(addr_width-1 downto 0) ;
    clk : in std_logic ;
    clken : in std_logic ;
    da : in std_logic_vector(data_width-1 downto 0) ;
    qa : out std_logic_vector(data_width-1 downto 0) ;
    qb : out std_logic_vector(data_width-1 downto 0) ;
    wea : in std_logic 
    
  );
  END COMPONENT;
END BLOCK_2R1W_RBW_pkg;
LIBRARY ieee;

  USE ieee.std_logic_1164.all;
  USE ieee.numeric_std.all;
ENTITY BLOCK_2R1W_RBW IS
  GENERIC (
    addr_width : integer := 8 ;
    data_width : integer := 7 ;
    depth : integer := 256 ;
    latency : integer := 1 
    
  );
  PORT (
    adra : in std_logic_vector(addr_width-1 downto 0) ;
    adrb : in std_logic_vector(addr_width-1 downto 0) ;
    clk : in std_logic ;
    clken : in std_logic ;
    da : in std_logic_vector(data_width-1 downto 0) ;
    qa : out std_logic_vector(data_width-1 downto 0) ;
    qb : out std_logic_vector(data_width-1 downto 0) ;
    wea : in std_logic 
    
  );
 END BLOCK_2R1W_RBW;
ARCHITECTURE rtl OF BLOCK_2R1W_RBW IS
  TYPE ram_t IS ARRAY (depth-1 DOWNTO 0) OF std_logic_vector(data_width-1 DOWNTO 0);
  SIGNAL mem : ram_t := (OTHERS => (OTHERS => '0'));
  ATTRIBUTE ram_style: STRING;
  ATTRIBUTE ram_style OF mem : SIGNAL IS "block";
  ATTRIBUTE syn_ramstyle: STRING;
  ATTRIBUTE syn_ramstyle OF mem : SIGNAL IS "block";
  
  SIGNAL ramqa : std_logic_vector(data_width-1 downto 0);
  SIGNAL ramqb : std_logic_vector(data_width-1 downto 0);
  
BEGIN
-- Port Map
-- rwA :: ADDRESS adra CLOCK clk ENABLE clken DATA_IN da DATA_OUT qa WRITE_ENABLE wea
-- readB :: ADDRESS adrb CLOCK clk ENABLE clken DATA_OUT qb

-- Access memory with non-registered inputs (latency = 1||2)
  IN_PIN :  IF latency < 3 GENERATE
  BEGIN
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
         IF (clken = '1') THEN
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (to_integer(unsigned(adra)) < depth) THEN
          --pragma translate_on
          ramqa <= mem(to_integer(unsigned(adra)));
          --pragma translate_off
          END IF;
          --pragma translate_on
          IF (wea = '1') THEN
            mem(to_integer(unsigned(adra))) <= da;
          END IF;
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (to_integer(unsigned(adrb)) < depth) THEN
          --pragma translate_on
          ramqb <= mem(to_integer(unsigned(adrb)));
          --pragma translate_off
          END IF;
          --pragma translate_on
        END IF;
      END IF;
    END PROCESS;
    
  END GENERATE IN_PIN; 

-- Register all non-clock inputs (latency = 3||4)
  IN_REG :  IF latency > 2 GENERATE
    SIGNAL adra_reg : std_logic_vector(addr_width-1 downto 0);
    SIGNAL da_reg : std_logic_vector(data_width-1 downto 0);
    SIGNAL wea_reg : std_logic;
    SIGNAL adrb_reg : std_logic_vector(addr_width-1 downto 0);
    
  BEGIN
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
        IF (clken = '1') THEN
          adra_reg <= adra;
          da_reg <= da;
          wea_reg <= wea;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
        IF (clken = '1') THEN
          adrb_reg <= adrb;
        END IF;
      END IF;
    END PROCESS;
    
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
         IF (clken = '1') THEN
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (to_integer(unsigned(adra_reg)) < depth) THEN
          --pragma translate_on
          ramqa <= mem(to_integer(unsigned(adra_reg)));
          --pragma translate_off
          END IF;
          --pragma translate_on
          IF (wea_reg = '1') THEN
            mem(to_integer(unsigned(adra_reg))) <= da_reg;
          END IF;
          -- workaround for simulation when read address out-of-range during inactive cycle
          --pragma translate_off
          IF (to_integer(unsigned(adrb_reg)) < depth) THEN
          --pragma translate_on
          ramqb <= mem(to_integer(unsigned(adrb_reg)));
          --pragma translate_off
          END IF;
          --pragma translate_on
        END IF;
      END IF;
    END PROCESS;
    
  END GENERATE IN_REG;

  out_ram : IF latency = 1 GENERATE
  BEGIN
    qa <= ramqa;
    qb <= ramqb;
    
  END GENERATE out_ram;

  out_reg1 : IF ((latency = 2) OR (latency = 3)) GENERATE
    SIGNAL tmpqa : std_logic_vector(data_width-1 downto 0);
    SIGNAL tmpqb : std_logic_vector(data_width-1 downto 0);
    
  BEGIN
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
        IF (clken = '1') THEN
          tmpqa <= ramqa;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
        IF (clken = '1') THEN
          tmpqb <= ramqb;
        END IF;
      END IF;
    END PROCESS;
    
    qa <= tmpqa;
    qb <= tmpqb;
    
  END GENERATE out_reg1;

  out_reg2 : IF latency = 4 GENERATE
    SIGNAL tmp1qa : std_logic_vector(data_width-1 downto 0);
    SIGNAL tmp1qb : std_logic_vector(data_width-1 downto 0);
    
    SIGNAL tmp2qa : std_logic_vector(data_width-1 downto 0);
    SIGNAL tmp2qb : std_logic_vector(data_width-1 downto 0);
    
  BEGIN
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
        IF (clken = '1') THEN
          tmp1qa <= ramqa;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
        IF (clken = '1') THEN
          tmp1qb <= ramqb;
        END IF;
      END IF;
    END PROCESS;
    
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
        IF (clken = '1') THEN
          tmp2qa <= tmp1qa;
        END IF;
      END IF;
    END PROCESS;
    PROCESS (clk)
    BEGIN
      IF (rising_edge(clk)) THEN
        IF (clken = '1') THEN
          tmp2qb <= tmp1qb;
        END IF;
      END IF;
    END PROCESS;
    
    qa <= tmp2qa;
    qb <= tmp2qb;
    
  END GENERATE out_reg2;


END rtl;

--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    10.5c/896140 Production Release
--  HLS Date:       Sun Sep  6 22:45:38 PDT 2020
-- 
--  Generated by:   jd4691@newnano.poly.edu
--  Generated date: Sun Sep 12 02:31:29 2021
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_134_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_134_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_134_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_134_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_133_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_133_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_133_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_133_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_132_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_132_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_132_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_132_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_131_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_131_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_131_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_131_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_130_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_130_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_130_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_130_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_129_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_129_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_129_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_129_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_128_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_128_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_128_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_128_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_127_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_127_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_127_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_127_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_126_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_126_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_126_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_126_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_125_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_125_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_125_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_125_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_124_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_124_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_124_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_124_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_123_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_123_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_123_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_123_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_122_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_122_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_122_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_122_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_121_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_121_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_121_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_121_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_120_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_120_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_120_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_120_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_119_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_119_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_119_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_119_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_118_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_118_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_118_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_118_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_117_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_117_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_117_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_117_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_116_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_116_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_116_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_116_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_115_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_115_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_115_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_115_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_114_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_114_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_114_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_114_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_113_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_113_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_113_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_113_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_112_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_112_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_112_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_112_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_111_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_111_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_111_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_111_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_110_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_110_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_110_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_110_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_109_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_109_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_109_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_109_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_108_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_108_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_108_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_108_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_107_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_107_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_107_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_107_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_106_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_106_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_106_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_106_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_105_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_105_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_105_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_105_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_104_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_104_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_104_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_104_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_103_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_103_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_103_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_103_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_102_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_102_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_102_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_102_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_101_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_101_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_101_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_101_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_100_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_100_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_100_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_100_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_99_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_99_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_99_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_99_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_98_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_98_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_98_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_98_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_97_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_97_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_97_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_97_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_96_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_96_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_96_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_96_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_95_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_95_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_95_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_95_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_94_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_94_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_94_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_94_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_93_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_93_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_93_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_93_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_92_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_92_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_92_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_92_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_91_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_91_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_91_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_91_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_90_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_90_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_90_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_90_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_89_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_89_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_89_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_89_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_88_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_88_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_88_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_88_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_87_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_87_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_87_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_87_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_86_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_86_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_86_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_86_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_85_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_85_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_85_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_85_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_84_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_84_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_84_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_84_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_83_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_83_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_83_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_83_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_82_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_82_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_82_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_82_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_81_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_81_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_81_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_81_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_80_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_80_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_80_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_80_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_79_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_79_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_79_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_79_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_78_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_78_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_78_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_78_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_77_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_77_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_77_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_77_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_76_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_76_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_76_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_76_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_75_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_75_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_75_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_75_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_74_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_74_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_74_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_74_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_73_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_73_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_73_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_73_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_72_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_72_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_72_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_72_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_71_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_71_4_32_16_16_32_1_gen IS
  PORT(
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_71_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_71_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_70_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_70_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_70_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_70_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_69_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_69_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_69_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_69_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_68_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_68_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_68_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_68_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_67_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_67_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_67_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_67_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_66_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_66_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_66_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_66_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_65_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_65_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_65_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_65_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_64_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_64_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_64_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_64_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_63_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_63_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_63_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_63_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_62_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_62_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_62_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_62_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_61_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_61_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_61_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_61_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_60_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_60_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_60_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_60_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_59_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_59_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_59_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_59_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_58_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_58_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_58_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_58_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_57_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_57_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_57_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_57_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_56_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_56_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_56_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_56_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_55_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_55_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_55_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_55_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_54_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_54_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_54_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_54_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_53_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_53_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_53_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_53_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_52_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_52_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_52_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_52_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_51_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_51_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_51_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_51_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_50_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_50_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_50_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_50_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_49_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_49_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_49_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_49_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_48_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_48_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_48_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_48_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_47_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_47_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_47_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_47_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_46_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_46_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_46_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_46_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_45_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_45_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_45_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_45_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_44_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_44_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_44_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_44_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_43_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_43_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_43_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_43_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_42_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_42_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_42_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_42_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_41_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_41_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_41_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_41_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_40_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_40_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_40_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_40_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_39_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_39_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_39_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_39_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_38_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_38_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_38_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_38_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_37_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_37_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_37_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_37_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_36_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_36_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_36_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_36_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_35_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_35_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_35_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_35_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_34_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_34_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_34_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_34_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_33_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_33_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_33_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_33_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_32_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_32_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_32_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_32_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_31_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_31_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_31_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_31_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_30_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_30_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_30_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_30_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_29_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_29_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_29_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_29_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_28_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_28_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_28_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_28_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_27_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_27_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_27_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_27_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_26_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_26_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_26_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_26_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_25_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_25_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_25_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_25_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_24_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_24_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_24_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_24_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_23_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_23_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_23_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_23_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_22_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_22_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_22_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_22_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_21_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_21_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_21_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_21_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_20_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_20_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_20_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_20_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_19_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_19_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_19_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_19_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_18_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_18_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_18_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_18_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_17_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_17_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_17_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_17_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_16_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_16_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_16_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_16_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_15_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_15_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_15_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_15_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_14_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_14_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_14_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_14_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_13_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_13_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_13_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_13_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_12_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_12_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_12_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_12_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_11_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_11_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_11_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_11_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_10_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_10_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_10_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_10_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_9_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_9_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_9_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_9_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_8_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_8_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_8_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_8_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_7_4_32_16_16_32_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_7_4_32_16_16_32_1_gen IS
  PORT(
    clken : OUT STD_LOGIC;
    qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea : OUT STD_LOGIC;
    da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    wea_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
    rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_7_4_32_16_16_32_1_gen;

ARCHITECTURE v29 OF peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_7_4_32_16_16_32_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  qa_d <= qa;
  wea <= (rwA_rw_ram_ir_internal_WMASK_B_d);
  da <= (da_d);
  adra <= (adra_d);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_core_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_core_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
    INNER_LOOP1_C_0_tr0 : IN STD_LOGIC;
    INNER_LOOP2_C_0_tr0 : IN STD_LOGIC;
    INNER_LOOP2_C_0_tr1 : IN STD_LOGIC;
    INNER_LOOP3_C_0_tr0 : IN STD_LOGIC;
    INNER_LOOP4_C_0_tr0 : IN STD_LOGIC;
    INNER_LOOP4_C_0_tr1 : IN STD_LOGIC
  );
END peaseNTT_core_core_fsm;

ARCHITECTURE v29 OF peaseNTT_core_core_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for peaseNTT_core_core_fsm_1
  TYPE peaseNTT_core_core_fsm_1_ST IS (main_C_0, STAGE_LOOP_C_0, INNER_LOOP1_C_0,
      STAGE_LOOP_C_1, INNER_LOOP2_C_0, STAGE_LOOP1_C_0, INNER_LOOP3_C_0, STAGE_LOOP1_C_1,
      INNER_LOOP4_C_0, main_C_1);

  SIGNAL state_var : peaseNTT_core_core_fsm_1_ST;
  SIGNAL state_var_NS : peaseNTT_core_core_fsm_1_ST;

BEGIN
  peaseNTT_core_core_fsm_1 : PROCESS (INNER_LOOP1_C_0_tr0, INNER_LOOP2_C_0_tr0, INNER_LOOP2_C_0_tr1,
      INNER_LOOP3_C_0_tr0, INNER_LOOP4_C_0_tr0, INNER_LOOP4_C_0_tr1, state_var)
  BEGIN
    CASE state_var IS
      WHEN STAGE_LOOP_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000010");
        state_var_NS <= INNER_LOOP1_C_0;
      WHEN INNER_LOOP1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000100");
        IF ( INNER_LOOP1_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP_C_1;
        ELSE
          state_var_NS <= INNER_LOOP1_C_0;
        END IF;
      WHEN STAGE_LOOP_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001000");
        state_var_NS <= INNER_LOOP2_C_0;
      WHEN INNER_LOOP2_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010000");
        IF ( INNER_LOOP2_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP1_C_0;
        ELSIF ( INNER_LOOP2_C_0_tr1 = '1' ) THEN
          state_var_NS <= INNER_LOOP2_C_0;
        ELSE
          state_var_NS <= STAGE_LOOP_C_0;
        END IF;
      WHEN STAGE_LOOP1_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100000");
        state_var_NS <= INNER_LOOP3_C_0;
      WHEN INNER_LOOP3_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000000");
        IF ( INNER_LOOP3_C_0_tr0 = '1' ) THEN
          state_var_NS <= STAGE_LOOP1_C_1;
        ELSE
          state_var_NS <= INNER_LOOP3_C_0;
        END IF;
      WHEN STAGE_LOOP1_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000000");
        state_var_NS <= INNER_LOOP4_C_0;
      WHEN INNER_LOOP4_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000000");
        IF ( INNER_LOOP4_C_0_tr0 = '1' ) THEN
          state_var_NS <= main_C_1;
        ELSIF ( INNER_LOOP4_C_0_tr1 = '1' ) THEN
          state_var_NS <= INNER_LOOP4_C_0;
        ELSE
          state_var_NS <= STAGE_LOOP1_C_0;
        END IF;
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000000");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000001");
        state_var_NS <= STAGE_LOOP_C_0;
    END CASE;
  END PROCESS peaseNTT_core_core_fsm_1;

  peaseNTT_core_core_fsm_1_REG : PROCESS (clk)
  BEGIN
    IF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        IF ( core_wen = '1' ) THEN
          state_var <= state_var_NS;
        END IF;
      END IF;
    END IF;
  END PROCESS peaseNTT_core_core_fsm_1_REG;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_staller
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_staller IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    core_wen : OUT STD_LOGIC;
    core_wten : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_1_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_2_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_3_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_4_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_5_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_6_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_7_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_8_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_9_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_10_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_11_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_12_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_13_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_14_i_wen_comp : IN STD_LOGIC;
    twiddle_rsc_0_15_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_8_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_9_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_10_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_11_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_12_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_13_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_14_i_wen_comp : IN STD_LOGIC;
    twiddle_h_rsc_0_15_i_wen_comp : IN STD_LOGIC
  );
END peaseNTT_core_staller;

ARCHITECTURE v29 OF peaseNTT_core_staller IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL core_wen_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL core_wten_reg : STD_LOGIC;

BEGIN
  -- Output Reader Assignments
  core_wen <= core_wen_drv;

  core_wen_drv <= twiddle_rsc_0_0_i_wen_comp AND twiddle_rsc_0_1_i_wen_comp AND twiddle_rsc_0_2_i_wen_comp
      AND twiddle_rsc_0_3_i_wen_comp AND twiddle_rsc_0_4_i_wen_comp AND twiddle_rsc_0_5_i_wen_comp
      AND twiddle_rsc_0_6_i_wen_comp AND twiddle_rsc_0_7_i_wen_comp AND twiddle_rsc_0_8_i_wen_comp
      AND twiddle_rsc_0_9_i_wen_comp AND twiddle_rsc_0_10_i_wen_comp AND twiddle_rsc_0_11_i_wen_comp
      AND twiddle_rsc_0_12_i_wen_comp AND twiddle_rsc_0_13_i_wen_comp AND twiddle_rsc_0_14_i_wen_comp
      AND twiddle_rsc_0_15_i_wen_comp AND twiddle_h_rsc_0_0_i_wen_comp AND twiddle_h_rsc_0_1_i_wen_comp
      AND twiddle_h_rsc_0_2_i_wen_comp AND twiddle_h_rsc_0_3_i_wen_comp AND twiddle_h_rsc_0_4_i_wen_comp
      AND twiddle_h_rsc_0_5_i_wen_comp AND twiddle_h_rsc_0_6_i_wen_comp AND twiddle_h_rsc_0_7_i_wen_comp
      AND twiddle_h_rsc_0_8_i_wen_comp AND twiddle_h_rsc_0_9_i_wen_comp AND twiddle_h_rsc_0_10_i_wen_comp
      AND twiddle_h_rsc_0_11_i_wen_comp AND twiddle_h_rsc_0_12_i_wen_comp AND twiddle_h_rsc_0_13_i_wen_comp
      AND twiddle_h_rsc_0_14_i_wen_comp AND twiddle_h_rsc_0_15_i_wen_comp;
  core_wten <= core_wten_reg;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        core_wten_reg <= '0';
      ELSE
        core_wten_reg <= NOT core_wen_drv;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_0_obj_twiddle_h_rsc_triosy_0_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_0_obj_twiddle_h_rsc_triosy_0_0_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_0_obj_twiddle_h_rsc_triosy_0_0_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_0_obj_twiddle_h_rsc_triosy_0_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_0_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_0_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_1_obj_twiddle_h_rsc_triosy_0_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_1_obj_twiddle_h_rsc_triosy_0_1_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_1_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_1_obj_twiddle_h_rsc_triosy_0_1_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_1_obj_twiddle_h_rsc_triosy_0_1_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_1_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_1_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_2_obj_twiddle_h_rsc_triosy_0_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_2_obj_twiddle_h_rsc_triosy_0_2_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_2_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_2_obj_twiddle_h_rsc_triosy_0_2_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_2_obj_twiddle_h_rsc_triosy_0_2_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_2_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_2_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_3_obj_twiddle_h_rsc_triosy_0_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_3_obj_twiddle_h_rsc_triosy_0_3_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_3_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_3_obj_twiddle_h_rsc_triosy_0_3_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_3_obj_twiddle_h_rsc_triosy_0_3_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_3_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_3_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_4_obj_twiddle_h_rsc_triosy_0_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_4_obj_twiddle_h_rsc_triosy_0_4_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_4_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_4_obj_twiddle_h_rsc_triosy_0_4_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_4_obj_twiddle_h_rsc_triosy_0_4_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_4_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_4_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_5_obj_twiddle_h_rsc_triosy_0_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_5_obj_twiddle_h_rsc_triosy_0_5_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_5_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_5_obj_twiddle_h_rsc_triosy_0_5_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_5_obj_twiddle_h_rsc_triosy_0_5_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_5_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_5_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_6_obj_twiddle_h_rsc_triosy_0_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_6_obj_twiddle_h_rsc_triosy_0_6_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_6_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_6_obj_twiddle_h_rsc_triosy_0_6_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_6_obj_twiddle_h_rsc_triosy_0_6_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_6_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_6_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_7_obj_twiddle_h_rsc_triosy_0_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_7_obj_twiddle_h_rsc_triosy_0_7_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_7_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_7_obj_twiddle_h_rsc_triosy_0_7_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_7_obj_twiddle_h_rsc_triosy_0_7_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_7_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_7_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_8_obj_twiddle_h_rsc_triosy_0_8_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_8_obj_twiddle_h_rsc_triosy_0_8_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_8_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_8_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_8_obj_twiddle_h_rsc_triosy_0_8_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_8_obj_twiddle_h_rsc_triosy_0_8_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_8_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_8_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_9_obj_twiddle_h_rsc_triosy_0_9_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_9_obj_twiddle_h_rsc_triosy_0_9_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_9_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_9_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_9_obj_twiddle_h_rsc_triosy_0_9_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_9_obj_twiddle_h_rsc_triosy_0_9_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_9_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_9_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_10_obj_twiddle_h_rsc_triosy_0_10_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_10_obj_twiddle_h_rsc_triosy_0_10_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_10_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_10_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_10_obj_twiddle_h_rsc_triosy_0_10_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_10_obj_twiddle_h_rsc_triosy_0_10_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_10_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_10_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_11_obj_twiddle_h_rsc_triosy_0_11_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_11_obj_twiddle_h_rsc_triosy_0_11_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_11_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_11_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_11_obj_twiddle_h_rsc_triosy_0_11_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_11_obj_twiddle_h_rsc_triosy_0_11_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_11_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_11_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_12_obj_twiddle_h_rsc_triosy_0_12_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_12_obj_twiddle_h_rsc_triosy_0_12_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_12_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_12_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_12_obj_twiddle_h_rsc_triosy_0_12_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_12_obj_twiddle_h_rsc_triosy_0_12_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_12_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_12_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_13_obj_twiddle_h_rsc_triosy_0_13_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_13_obj_twiddle_h_rsc_triosy_0_13_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_13_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_13_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_13_obj_twiddle_h_rsc_triosy_0_13_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_13_obj_twiddle_h_rsc_triosy_0_13_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_13_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_13_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_14_obj_twiddle_h_rsc_triosy_0_14_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_14_obj_twiddle_h_rsc_triosy_0_14_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_14_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_14_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_14_obj_twiddle_h_rsc_triosy_0_14_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_14_obj_twiddle_h_rsc_triosy_0_14_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_14_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_14_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_15_obj_twiddle_h_rsc_triosy_0_15_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_15_obj_twiddle_h_rsc_triosy_0_15_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_15_obj_iswt0 : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_15_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_15_obj_twiddle_h_rsc_triosy_0_15_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_15_obj_twiddle_h_rsc_triosy_0_15_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_h_rsc_triosy_0_15_obj_ld_core_sct <= twiddle_h_rsc_triosy_0_15_obj_iswt0
      AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_0_obj_twiddle_rsc_triosy_0_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_0_obj_twiddle_rsc_triosy_0_0_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_0_obj_twiddle_rsc_triosy_0_0_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_0_obj_twiddle_rsc_triosy_0_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_0_obj_ld_core_sct <= twiddle_rsc_triosy_0_0_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_1_obj_twiddle_rsc_triosy_0_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_1_obj_twiddle_rsc_triosy_0_1_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_1_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_1_obj_twiddle_rsc_triosy_0_1_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_1_obj_twiddle_rsc_triosy_0_1_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_1_obj_ld_core_sct <= twiddle_rsc_triosy_0_1_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_2_obj_twiddle_rsc_triosy_0_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_2_obj_twiddle_rsc_triosy_0_2_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_2_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_2_obj_twiddle_rsc_triosy_0_2_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_2_obj_twiddle_rsc_triosy_0_2_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_2_obj_ld_core_sct <= twiddle_rsc_triosy_0_2_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_3_obj_twiddle_rsc_triosy_0_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_3_obj_twiddle_rsc_triosy_0_3_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_3_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_3_obj_twiddle_rsc_triosy_0_3_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_3_obj_twiddle_rsc_triosy_0_3_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_3_obj_ld_core_sct <= twiddle_rsc_triosy_0_3_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_4_obj_twiddle_rsc_triosy_0_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_4_obj_twiddle_rsc_triosy_0_4_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_4_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_4_obj_twiddle_rsc_triosy_0_4_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_4_obj_twiddle_rsc_triosy_0_4_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_4_obj_ld_core_sct <= twiddle_rsc_triosy_0_4_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_5_obj_twiddle_rsc_triosy_0_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_5_obj_twiddle_rsc_triosy_0_5_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_5_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_5_obj_twiddle_rsc_triosy_0_5_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_5_obj_twiddle_rsc_triosy_0_5_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_5_obj_ld_core_sct <= twiddle_rsc_triosy_0_5_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_6_obj_twiddle_rsc_triosy_0_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_6_obj_twiddle_rsc_triosy_0_6_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_6_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_6_obj_twiddle_rsc_triosy_0_6_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_6_obj_twiddle_rsc_triosy_0_6_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_6_obj_ld_core_sct <= twiddle_rsc_triosy_0_6_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_7_obj_twiddle_rsc_triosy_0_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_7_obj_twiddle_rsc_triosy_0_7_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_7_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_7_obj_twiddle_rsc_triosy_0_7_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_7_obj_twiddle_rsc_triosy_0_7_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_7_obj_ld_core_sct <= twiddle_rsc_triosy_0_7_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_8_obj_twiddle_rsc_triosy_0_8_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_8_obj_twiddle_rsc_triosy_0_8_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_8_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_8_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_8_obj_twiddle_rsc_triosy_0_8_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_8_obj_twiddle_rsc_triosy_0_8_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_8_obj_ld_core_sct <= twiddle_rsc_triosy_0_8_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_9_obj_twiddle_rsc_triosy_0_9_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_9_obj_twiddle_rsc_triosy_0_9_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_9_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_9_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_9_obj_twiddle_rsc_triosy_0_9_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_9_obj_twiddle_rsc_triosy_0_9_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_9_obj_ld_core_sct <= twiddle_rsc_triosy_0_9_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_10_obj_twiddle_rsc_triosy_0_10_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_10_obj_twiddle_rsc_triosy_0_10_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_10_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_10_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_10_obj_twiddle_rsc_triosy_0_10_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_10_obj_twiddle_rsc_triosy_0_10_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_10_obj_ld_core_sct <= twiddle_rsc_triosy_0_10_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_11_obj_twiddle_rsc_triosy_0_11_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_11_obj_twiddle_rsc_triosy_0_11_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_11_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_11_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_11_obj_twiddle_rsc_triosy_0_11_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_11_obj_twiddle_rsc_triosy_0_11_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_11_obj_ld_core_sct <= twiddle_rsc_triosy_0_11_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_12_obj_twiddle_rsc_triosy_0_12_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_12_obj_twiddle_rsc_triosy_0_12_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_12_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_12_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_12_obj_twiddle_rsc_triosy_0_12_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_12_obj_twiddle_rsc_triosy_0_12_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_12_obj_ld_core_sct <= twiddle_rsc_triosy_0_12_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_13_obj_twiddle_rsc_triosy_0_13_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_13_obj_twiddle_rsc_triosy_0_13_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_13_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_13_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_13_obj_twiddle_rsc_triosy_0_13_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_13_obj_twiddle_rsc_triosy_0_13_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_13_obj_ld_core_sct <= twiddle_rsc_triosy_0_13_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_14_obj_twiddle_rsc_triosy_0_14_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_14_obj_twiddle_rsc_triosy_0_14_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_14_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_14_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_14_obj_twiddle_rsc_triosy_0_14_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_14_obj_twiddle_rsc_triosy_0_14_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_14_obj_ld_core_sct <= twiddle_rsc_triosy_0_14_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_15_obj_twiddle_rsc_triosy_0_15_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_15_obj_twiddle_rsc_triosy_0_15_wait_ctrl
    IS
  PORT(
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_15_obj_iswt0 : IN STD_LOGIC;
    twiddle_rsc_triosy_0_15_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_15_obj_twiddle_rsc_triosy_0_15_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_15_obj_twiddle_rsc_triosy_0_15_wait_ctrl
    IS
  -- Default Constants

BEGIN
  twiddle_rsc_triosy_0_15_obj_ld_core_sct <= twiddle_rsc_triosy_0_15_obj_iswt0 AND
      (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_r_rsc_triosy_obj_r_rsc_triosy_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_r_rsc_triosy_obj_r_rsc_triosy_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    r_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
    r_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_r_rsc_triosy_obj_r_rsc_triosy_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_r_rsc_triosy_obj_r_rsc_triosy_wait_ctrl IS
  -- Default Constants

BEGIN
  r_rsc_triosy_obj_ld_core_sct <= r_rsc_triosy_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_p_rsc_triosy_obj_p_rsc_triosy_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_p_rsc_triosy_obj_p_rsc_triosy_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    p_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
    p_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_p_rsc_triosy_obj_p_rsc_triosy_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_p_rsc_triosy_obj_p_rsc_triosy_wait_ctrl IS
  -- Default Constants

BEGIN
  p_rsc_triosy_obj_ld_core_sct <= p_rsc_triosy_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_0_obj_xt_rsc_triosy_0_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_0_obj_xt_rsc_triosy_0_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_0_obj_xt_rsc_triosy_0_0_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_0_obj_xt_rsc_triosy_0_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_0_obj_ld_core_sct <= xt_rsc_triosy_0_0_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_1_obj_xt_rsc_triosy_0_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_1_obj_xt_rsc_triosy_0_1_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_1_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_1_obj_xt_rsc_triosy_0_1_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_1_obj_xt_rsc_triosy_0_1_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_1_obj_ld_core_sct <= xt_rsc_triosy_0_1_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_2_obj_xt_rsc_triosy_0_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_2_obj_xt_rsc_triosy_0_2_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_2_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_2_obj_xt_rsc_triosy_0_2_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_2_obj_xt_rsc_triosy_0_2_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_2_obj_ld_core_sct <= xt_rsc_triosy_0_2_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_3_obj_xt_rsc_triosy_0_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_3_obj_xt_rsc_triosy_0_3_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_3_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_3_obj_xt_rsc_triosy_0_3_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_3_obj_xt_rsc_triosy_0_3_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_3_obj_ld_core_sct <= xt_rsc_triosy_0_3_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_4_obj_xt_rsc_triosy_0_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_4_obj_xt_rsc_triosy_0_4_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_4_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_4_obj_xt_rsc_triosy_0_4_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_4_obj_xt_rsc_triosy_0_4_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_4_obj_ld_core_sct <= xt_rsc_triosy_0_4_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_5_obj_xt_rsc_triosy_0_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_5_obj_xt_rsc_triosy_0_5_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_5_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_5_obj_xt_rsc_triosy_0_5_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_5_obj_xt_rsc_triosy_0_5_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_5_obj_ld_core_sct <= xt_rsc_triosy_0_5_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_6_obj_xt_rsc_triosy_0_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_6_obj_xt_rsc_triosy_0_6_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_6_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_6_obj_xt_rsc_triosy_0_6_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_6_obj_xt_rsc_triosy_0_6_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_6_obj_ld_core_sct <= xt_rsc_triosy_0_6_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_7_obj_xt_rsc_triosy_0_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_7_obj_xt_rsc_triosy_0_7_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_7_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_7_obj_xt_rsc_triosy_0_7_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_7_obj_xt_rsc_triosy_0_7_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_7_obj_ld_core_sct <= xt_rsc_triosy_0_7_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_8_obj_xt_rsc_triosy_0_8_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_8_obj_xt_rsc_triosy_0_8_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_8_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_8_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_8_obj_xt_rsc_triosy_0_8_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_8_obj_xt_rsc_triosy_0_8_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_8_obj_ld_core_sct <= xt_rsc_triosy_0_8_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_9_obj_xt_rsc_triosy_0_9_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_9_obj_xt_rsc_triosy_0_9_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_9_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_9_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_9_obj_xt_rsc_triosy_0_9_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_9_obj_xt_rsc_triosy_0_9_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_9_obj_ld_core_sct <= xt_rsc_triosy_0_9_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_10_obj_xt_rsc_triosy_0_10_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_10_obj_xt_rsc_triosy_0_10_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_10_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_10_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_10_obj_xt_rsc_triosy_0_10_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_10_obj_xt_rsc_triosy_0_10_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_10_obj_ld_core_sct <= xt_rsc_triosy_0_10_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_11_obj_xt_rsc_triosy_0_11_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_11_obj_xt_rsc_triosy_0_11_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_11_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_11_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_11_obj_xt_rsc_triosy_0_11_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_11_obj_xt_rsc_triosy_0_11_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_11_obj_ld_core_sct <= xt_rsc_triosy_0_11_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_12_obj_xt_rsc_triosy_0_12_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_12_obj_xt_rsc_triosy_0_12_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_12_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_12_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_12_obj_xt_rsc_triosy_0_12_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_12_obj_xt_rsc_triosy_0_12_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_12_obj_ld_core_sct <= xt_rsc_triosy_0_12_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_13_obj_xt_rsc_triosy_0_13_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_13_obj_xt_rsc_triosy_0_13_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_13_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_13_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_13_obj_xt_rsc_triosy_0_13_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_13_obj_xt_rsc_triosy_0_13_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_13_obj_ld_core_sct <= xt_rsc_triosy_0_13_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_14_obj_xt_rsc_triosy_0_14_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_14_obj_xt_rsc_triosy_0_14_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_14_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_14_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_14_obj_xt_rsc_triosy_0_14_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_14_obj_xt_rsc_triosy_0_14_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_14_obj_ld_core_sct <= xt_rsc_triosy_0_14_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_15_obj_xt_rsc_triosy_0_15_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_15_obj_xt_rsc_triosy_0_15_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_15_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_15_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_15_obj_xt_rsc_triosy_0_15_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_15_obj_xt_rsc_triosy_0_15_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_15_obj_ld_core_sct <= xt_rsc_triosy_0_15_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_16_obj_xt_rsc_triosy_0_16_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_16_obj_xt_rsc_triosy_0_16_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_16_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_16_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_16_obj_xt_rsc_triosy_0_16_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_16_obj_xt_rsc_triosy_0_16_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_16_obj_ld_core_sct <= xt_rsc_triosy_0_16_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_17_obj_xt_rsc_triosy_0_17_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_17_obj_xt_rsc_triosy_0_17_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_17_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_17_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_17_obj_xt_rsc_triosy_0_17_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_17_obj_xt_rsc_triosy_0_17_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_17_obj_ld_core_sct <= xt_rsc_triosy_0_17_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_18_obj_xt_rsc_triosy_0_18_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_18_obj_xt_rsc_triosy_0_18_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_18_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_18_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_18_obj_xt_rsc_triosy_0_18_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_18_obj_xt_rsc_triosy_0_18_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_18_obj_ld_core_sct <= xt_rsc_triosy_0_18_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_19_obj_xt_rsc_triosy_0_19_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_19_obj_xt_rsc_triosy_0_19_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_19_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_19_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_19_obj_xt_rsc_triosy_0_19_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_19_obj_xt_rsc_triosy_0_19_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_19_obj_ld_core_sct <= xt_rsc_triosy_0_19_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_20_obj_xt_rsc_triosy_0_20_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_20_obj_xt_rsc_triosy_0_20_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_20_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_20_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_20_obj_xt_rsc_triosy_0_20_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_20_obj_xt_rsc_triosy_0_20_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_20_obj_ld_core_sct <= xt_rsc_triosy_0_20_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_21_obj_xt_rsc_triosy_0_21_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_21_obj_xt_rsc_triosy_0_21_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_21_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_21_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_21_obj_xt_rsc_triosy_0_21_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_21_obj_xt_rsc_triosy_0_21_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_21_obj_ld_core_sct <= xt_rsc_triosy_0_21_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_22_obj_xt_rsc_triosy_0_22_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_22_obj_xt_rsc_triosy_0_22_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_22_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_22_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_22_obj_xt_rsc_triosy_0_22_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_22_obj_xt_rsc_triosy_0_22_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_22_obj_ld_core_sct <= xt_rsc_triosy_0_22_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_23_obj_xt_rsc_triosy_0_23_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_23_obj_xt_rsc_triosy_0_23_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_23_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_23_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_23_obj_xt_rsc_triosy_0_23_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_23_obj_xt_rsc_triosy_0_23_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_23_obj_ld_core_sct <= xt_rsc_triosy_0_23_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_24_obj_xt_rsc_triosy_0_24_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_24_obj_xt_rsc_triosy_0_24_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_24_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_24_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_24_obj_xt_rsc_triosy_0_24_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_24_obj_xt_rsc_triosy_0_24_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_24_obj_ld_core_sct <= xt_rsc_triosy_0_24_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_25_obj_xt_rsc_triosy_0_25_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_25_obj_xt_rsc_triosy_0_25_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_25_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_25_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_25_obj_xt_rsc_triosy_0_25_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_25_obj_xt_rsc_triosy_0_25_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_25_obj_ld_core_sct <= xt_rsc_triosy_0_25_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_26_obj_xt_rsc_triosy_0_26_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_26_obj_xt_rsc_triosy_0_26_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_26_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_26_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_26_obj_xt_rsc_triosy_0_26_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_26_obj_xt_rsc_triosy_0_26_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_26_obj_ld_core_sct <= xt_rsc_triosy_0_26_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_27_obj_xt_rsc_triosy_0_27_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_27_obj_xt_rsc_triosy_0_27_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_27_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_27_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_27_obj_xt_rsc_triosy_0_27_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_27_obj_xt_rsc_triosy_0_27_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_27_obj_ld_core_sct <= xt_rsc_triosy_0_27_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_28_obj_xt_rsc_triosy_0_28_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_28_obj_xt_rsc_triosy_0_28_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_28_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_28_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_28_obj_xt_rsc_triosy_0_28_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_28_obj_xt_rsc_triosy_0_28_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_28_obj_ld_core_sct <= xt_rsc_triosy_0_28_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_29_obj_xt_rsc_triosy_0_29_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_29_obj_xt_rsc_triosy_0_29_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_29_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_29_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_29_obj_xt_rsc_triosy_0_29_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_29_obj_xt_rsc_triosy_0_29_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_29_obj_ld_core_sct <= xt_rsc_triosy_0_29_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_30_obj_xt_rsc_triosy_0_30_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_30_obj_xt_rsc_triosy_0_30_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_30_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_30_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_30_obj_xt_rsc_triosy_0_30_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_30_obj_xt_rsc_triosy_0_30_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_30_obj_ld_core_sct <= xt_rsc_triosy_0_30_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_31_obj_xt_rsc_triosy_0_31_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_31_obj_xt_rsc_triosy_0_31_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_31_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_0_31_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_31_obj_xt_rsc_triosy_0_31_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_31_obj_xt_rsc_triosy_0_31_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_0_31_obj_ld_core_sct <= xt_rsc_triosy_0_31_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_0_obj_xt_rsc_triosy_1_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_0_obj_xt_rsc_triosy_1_0_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_0_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_0_obj_xt_rsc_triosy_1_0_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_0_obj_xt_rsc_triosy_1_0_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_0_obj_ld_core_sct <= xt_rsc_triosy_1_0_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_1_obj_xt_rsc_triosy_1_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_1_obj_xt_rsc_triosy_1_1_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_1_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_1_obj_xt_rsc_triosy_1_1_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_1_obj_xt_rsc_triosy_1_1_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_1_obj_ld_core_sct <= xt_rsc_triosy_1_1_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_2_obj_xt_rsc_triosy_1_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_2_obj_xt_rsc_triosy_1_2_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_2_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_2_obj_xt_rsc_triosy_1_2_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_2_obj_xt_rsc_triosy_1_2_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_2_obj_ld_core_sct <= xt_rsc_triosy_1_2_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_3_obj_xt_rsc_triosy_1_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_3_obj_xt_rsc_triosy_1_3_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_3_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_3_obj_xt_rsc_triosy_1_3_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_3_obj_xt_rsc_triosy_1_3_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_3_obj_ld_core_sct <= xt_rsc_triosy_1_3_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_4_obj_xt_rsc_triosy_1_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_4_obj_xt_rsc_triosy_1_4_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_4_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_4_obj_xt_rsc_triosy_1_4_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_4_obj_xt_rsc_triosy_1_4_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_4_obj_ld_core_sct <= xt_rsc_triosy_1_4_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_5_obj_xt_rsc_triosy_1_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_5_obj_xt_rsc_triosy_1_5_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_5_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_5_obj_xt_rsc_triosy_1_5_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_5_obj_xt_rsc_triosy_1_5_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_5_obj_ld_core_sct <= xt_rsc_triosy_1_5_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_6_obj_xt_rsc_triosy_1_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_6_obj_xt_rsc_triosy_1_6_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_6_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_6_obj_xt_rsc_triosy_1_6_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_6_obj_xt_rsc_triosy_1_6_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_6_obj_ld_core_sct <= xt_rsc_triosy_1_6_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_7_obj_xt_rsc_triosy_1_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_7_obj_xt_rsc_triosy_1_7_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_7_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_7_obj_xt_rsc_triosy_1_7_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_7_obj_xt_rsc_triosy_1_7_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_7_obj_ld_core_sct <= xt_rsc_triosy_1_7_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_8_obj_xt_rsc_triosy_1_8_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_8_obj_xt_rsc_triosy_1_8_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_8_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_8_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_8_obj_xt_rsc_triosy_1_8_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_8_obj_xt_rsc_triosy_1_8_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_8_obj_ld_core_sct <= xt_rsc_triosy_1_8_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_9_obj_xt_rsc_triosy_1_9_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_9_obj_xt_rsc_triosy_1_9_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_9_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_9_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_9_obj_xt_rsc_triosy_1_9_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_9_obj_xt_rsc_triosy_1_9_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_9_obj_ld_core_sct <= xt_rsc_triosy_1_9_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_10_obj_xt_rsc_triosy_1_10_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_10_obj_xt_rsc_triosy_1_10_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_10_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_10_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_10_obj_xt_rsc_triosy_1_10_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_10_obj_xt_rsc_triosy_1_10_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_10_obj_ld_core_sct <= xt_rsc_triosy_1_10_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_11_obj_xt_rsc_triosy_1_11_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_11_obj_xt_rsc_triosy_1_11_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_11_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_11_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_11_obj_xt_rsc_triosy_1_11_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_11_obj_xt_rsc_triosy_1_11_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_11_obj_ld_core_sct <= xt_rsc_triosy_1_11_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_12_obj_xt_rsc_triosy_1_12_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_12_obj_xt_rsc_triosy_1_12_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_12_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_12_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_12_obj_xt_rsc_triosy_1_12_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_12_obj_xt_rsc_triosy_1_12_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_12_obj_ld_core_sct <= xt_rsc_triosy_1_12_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_13_obj_xt_rsc_triosy_1_13_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_13_obj_xt_rsc_triosy_1_13_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_13_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_13_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_13_obj_xt_rsc_triosy_1_13_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_13_obj_xt_rsc_triosy_1_13_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_13_obj_ld_core_sct <= xt_rsc_triosy_1_13_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_14_obj_xt_rsc_triosy_1_14_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_14_obj_xt_rsc_triosy_1_14_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_14_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_14_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_14_obj_xt_rsc_triosy_1_14_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_14_obj_xt_rsc_triosy_1_14_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_14_obj_ld_core_sct <= xt_rsc_triosy_1_14_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_15_obj_xt_rsc_triosy_1_15_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_15_obj_xt_rsc_triosy_1_15_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_15_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_15_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_15_obj_xt_rsc_triosy_1_15_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_15_obj_xt_rsc_triosy_1_15_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_15_obj_ld_core_sct <= xt_rsc_triosy_1_15_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_16_obj_xt_rsc_triosy_1_16_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_16_obj_xt_rsc_triosy_1_16_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_16_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_16_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_16_obj_xt_rsc_triosy_1_16_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_16_obj_xt_rsc_triosy_1_16_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_16_obj_ld_core_sct <= xt_rsc_triosy_1_16_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_17_obj_xt_rsc_triosy_1_17_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_17_obj_xt_rsc_triosy_1_17_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_17_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_17_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_17_obj_xt_rsc_triosy_1_17_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_17_obj_xt_rsc_triosy_1_17_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_17_obj_ld_core_sct <= xt_rsc_triosy_1_17_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_18_obj_xt_rsc_triosy_1_18_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_18_obj_xt_rsc_triosy_1_18_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_18_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_18_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_18_obj_xt_rsc_triosy_1_18_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_18_obj_xt_rsc_triosy_1_18_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_18_obj_ld_core_sct <= xt_rsc_triosy_1_18_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_19_obj_xt_rsc_triosy_1_19_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_19_obj_xt_rsc_triosy_1_19_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_19_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_19_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_19_obj_xt_rsc_triosy_1_19_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_19_obj_xt_rsc_triosy_1_19_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_19_obj_ld_core_sct <= xt_rsc_triosy_1_19_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_20_obj_xt_rsc_triosy_1_20_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_20_obj_xt_rsc_triosy_1_20_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_20_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_20_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_20_obj_xt_rsc_triosy_1_20_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_20_obj_xt_rsc_triosy_1_20_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_20_obj_ld_core_sct <= xt_rsc_triosy_1_20_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_21_obj_xt_rsc_triosy_1_21_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_21_obj_xt_rsc_triosy_1_21_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_21_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_21_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_21_obj_xt_rsc_triosy_1_21_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_21_obj_xt_rsc_triosy_1_21_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_21_obj_ld_core_sct <= xt_rsc_triosy_1_21_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_22_obj_xt_rsc_triosy_1_22_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_22_obj_xt_rsc_triosy_1_22_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_22_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_22_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_22_obj_xt_rsc_triosy_1_22_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_22_obj_xt_rsc_triosy_1_22_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_22_obj_ld_core_sct <= xt_rsc_triosy_1_22_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_23_obj_xt_rsc_triosy_1_23_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_23_obj_xt_rsc_triosy_1_23_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_23_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_23_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_23_obj_xt_rsc_triosy_1_23_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_23_obj_xt_rsc_triosy_1_23_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_23_obj_ld_core_sct <= xt_rsc_triosy_1_23_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_24_obj_xt_rsc_triosy_1_24_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_24_obj_xt_rsc_triosy_1_24_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_24_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_24_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_24_obj_xt_rsc_triosy_1_24_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_24_obj_xt_rsc_triosy_1_24_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_24_obj_ld_core_sct <= xt_rsc_triosy_1_24_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_25_obj_xt_rsc_triosy_1_25_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_25_obj_xt_rsc_triosy_1_25_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_25_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_25_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_25_obj_xt_rsc_triosy_1_25_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_25_obj_xt_rsc_triosy_1_25_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_25_obj_ld_core_sct <= xt_rsc_triosy_1_25_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_26_obj_xt_rsc_triosy_1_26_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_26_obj_xt_rsc_triosy_1_26_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_26_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_26_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_26_obj_xt_rsc_triosy_1_26_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_26_obj_xt_rsc_triosy_1_26_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_26_obj_ld_core_sct <= xt_rsc_triosy_1_26_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_27_obj_xt_rsc_triosy_1_27_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_27_obj_xt_rsc_triosy_1_27_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_27_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_27_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_27_obj_xt_rsc_triosy_1_27_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_27_obj_xt_rsc_triosy_1_27_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_27_obj_ld_core_sct <= xt_rsc_triosy_1_27_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_28_obj_xt_rsc_triosy_1_28_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_28_obj_xt_rsc_triosy_1_28_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_28_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_28_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_28_obj_xt_rsc_triosy_1_28_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_28_obj_xt_rsc_triosy_1_28_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_28_obj_ld_core_sct <= xt_rsc_triosy_1_28_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_29_obj_xt_rsc_triosy_1_29_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_29_obj_xt_rsc_triosy_1_29_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_29_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_29_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_29_obj_xt_rsc_triosy_1_29_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_29_obj_xt_rsc_triosy_1_29_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_29_obj_ld_core_sct <= xt_rsc_triosy_1_29_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_30_obj_xt_rsc_triosy_1_30_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_30_obj_xt_rsc_triosy_1_30_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_30_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_30_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_30_obj_xt_rsc_triosy_1_30_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_30_obj_xt_rsc_triosy_1_30_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_30_obj_ld_core_sct <= xt_rsc_triosy_1_30_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_31_obj_xt_rsc_triosy_1_31_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_31_obj_xt_rsc_triosy_1_31_wait_ctrl IS
  PORT(
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_31_obj_iswt0 : IN STD_LOGIC;
    xt_rsc_triosy_1_31_obj_ld_core_sct : OUT STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_31_obj_xt_rsc_triosy_1_31_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_31_obj_xt_rsc_triosy_1_31_wait_ctrl
    IS
  -- Default Constants

BEGIN
  xt_rsc_triosy_1_31_obj_ld_core_sct <= xt_rsc_triosy_1_31_obj_iswt0 AND (NOT core_wten);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_15_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_15_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_15_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_15_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_15_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_15_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_15_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_15_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp
    IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_15_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_15_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_15_tw_h_butterFly2_15_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_15_i_bcwt <= twiddle_h_rsc_0_15_i_bcwt_drv;

  twiddle_h_rsc_0_15_i_wen_comp <= (NOT twiddle_h_rsc_0_15_i_oswt) OR twiddle_h_rsc_0_15_i_biwt
      OR twiddle_h_rsc_0_15_i_bcwt_drv;
  butterFly2_15_tw_h_butterFly2_15_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_15_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_15_i_s_raddr_core_sct);
  twiddle_h_rsc_0_15_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_15_tw_h_butterFly2_15_tw_h_and_nl));
  twiddle_h_rsc_0_15_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_15_i_s_din, twiddle_h_rsc_0_15_i_s_din_bfwt,
      twiddle_h_rsc_0_15_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_15_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_15_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_15_i_bcwt_drv OR
            twiddle_h_rsc_0_15_i_biwt)) OR twiddle_h_rsc_0_15_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_15_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_15_i_s_din_bfwt <= twiddle_h_rsc_0_15_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_15_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_15_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_15_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_15_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_15_i_bdwt <= twiddle_h_rsc_0_15_i_oswt AND core_wen;
  twiddle_h_rsc_0_15_i_biwt <= twiddle_h_rsc_0_15_i_ogwt AND twiddle_h_rsc_0_15_i_s_rrdy;
  twiddle_h_rsc_0_15_i_ogwt <= twiddle_h_rsc_0_15_i_oswt AND (NOT twiddle_h_rsc_0_15_i_bcwt);
  twiddle_h_rsc_0_15_i_s_re_core_sct <= twiddle_h_rsc_0_15_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_14_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_14_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_14_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_14_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_14_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_14_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_14_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_14_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp
    IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_14_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_14_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_14_tw_h_butterFly2_14_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_14_i_bcwt <= twiddle_h_rsc_0_14_i_bcwt_drv;

  twiddle_h_rsc_0_14_i_wen_comp <= (NOT twiddle_h_rsc_0_14_i_oswt) OR twiddle_h_rsc_0_14_i_biwt
      OR twiddle_h_rsc_0_14_i_bcwt_drv;
  butterFly2_14_tw_h_butterFly2_14_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_14_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_14_i_s_raddr_core_sct);
  twiddle_h_rsc_0_14_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_14_tw_h_butterFly2_14_tw_h_and_nl));
  twiddle_h_rsc_0_14_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_14_i_s_din, twiddle_h_rsc_0_14_i_s_din_bfwt,
      twiddle_h_rsc_0_14_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_14_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_14_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_14_i_bcwt_drv OR
            twiddle_h_rsc_0_14_i_biwt)) OR twiddle_h_rsc_0_14_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_14_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_14_i_s_din_bfwt <= twiddle_h_rsc_0_14_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_14_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_14_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_14_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_14_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_14_i_bdwt <= twiddle_h_rsc_0_14_i_oswt AND core_wen;
  twiddle_h_rsc_0_14_i_biwt <= twiddle_h_rsc_0_14_i_ogwt AND twiddle_h_rsc_0_14_i_s_rrdy;
  twiddle_h_rsc_0_14_i_ogwt <= twiddle_h_rsc_0_14_i_oswt AND (NOT twiddle_h_rsc_0_14_i_bcwt);
  twiddle_h_rsc_0_14_i_s_re_core_sct <= twiddle_h_rsc_0_14_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_13_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_13_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_13_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_13_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_13_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_13_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_13_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_13_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp
    IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_13_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_13_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_13_tw_h_butterFly2_13_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_13_i_bcwt <= twiddle_h_rsc_0_13_i_bcwt_drv;

  twiddle_h_rsc_0_13_i_wen_comp <= (NOT twiddle_h_rsc_0_13_i_oswt) OR twiddle_h_rsc_0_13_i_biwt
      OR twiddle_h_rsc_0_13_i_bcwt_drv;
  butterFly2_13_tw_h_butterFly2_13_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_13_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_13_i_s_raddr_core_sct);
  twiddle_h_rsc_0_13_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_13_tw_h_butterFly2_13_tw_h_and_nl));
  twiddle_h_rsc_0_13_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_13_i_s_din, twiddle_h_rsc_0_13_i_s_din_bfwt,
      twiddle_h_rsc_0_13_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_13_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_13_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_13_i_bcwt_drv OR
            twiddle_h_rsc_0_13_i_biwt)) OR twiddle_h_rsc_0_13_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_13_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_13_i_s_din_bfwt <= twiddle_h_rsc_0_13_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_13_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_13_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_13_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_13_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_13_i_bdwt <= twiddle_h_rsc_0_13_i_oswt AND core_wen;
  twiddle_h_rsc_0_13_i_biwt <= twiddle_h_rsc_0_13_i_ogwt AND twiddle_h_rsc_0_13_i_s_rrdy;
  twiddle_h_rsc_0_13_i_ogwt <= twiddle_h_rsc_0_13_i_oswt AND (NOT twiddle_h_rsc_0_13_i_bcwt);
  twiddle_h_rsc_0_13_i_s_re_core_sct <= twiddle_h_rsc_0_13_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_12_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_12_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_12_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_12_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_12_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_12_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_12_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_12_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp
    IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_12_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_12_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_12_tw_h_butterFly2_12_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_12_i_bcwt <= twiddle_h_rsc_0_12_i_bcwt_drv;

  twiddle_h_rsc_0_12_i_wen_comp <= (NOT twiddle_h_rsc_0_12_i_oswt) OR twiddle_h_rsc_0_12_i_biwt
      OR twiddle_h_rsc_0_12_i_bcwt_drv;
  butterFly2_12_tw_h_butterFly2_12_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_12_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_12_i_s_raddr_core_sct);
  twiddle_h_rsc_0_12_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_12_tw_h_butterFly2_12_tw_h_and_nl));
  twiddle_h_rsc_0_12_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_12_i_s_din, twiddle_h_rsc_0_12_i_s_din_bfwt,
      twiddle_h_rsc_0_12_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_12_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_12_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_12_i_bcwt_drv OR
            twiddle_h_rsc_0_12_i_biwt)) OR twiddle_h_rsc_0_12_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_12_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_12_i_s_din_bfwt <= twiddle_h_rsc_0_12_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_12_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_12_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_12_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_12_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_12_i_bdwt <= twiddle_h_rsc_0_12_i_oswt AND core_wen;
  twiddle_h_rsc_0_12_i_biwt <= twiddle_h_rsc_0_12_i_ogwt AND twiddle_h_rsc_0_12_i_s_rrdy;
  twiddle_h_rsc_0_12_i_ogwt <= twiddle_h_rsc_0_12_i_oswt AND (NOT twiddle_h_rsc_0_12_i_bcwt);
  twiddle_h_rsc_0_12_i_s_re_core_sct <= twiddle_h_rsc_0_12_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_11_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_11_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_11_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_11_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_11_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_11_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_11_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_11_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp
    IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_11_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_11_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_11_tw_h_butterFly2_11_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_11_i_bcwt <= twiddle_h_rsc_0_11_i_bcwt_drv;

  twiddle_h_rsc_0_11_i_wen_comp <= (NOT twiddle_h_rsc_0_11_i_oswt) OR twiddle_h_rsc_0_11_i_biwt
      OR twiddle_h_rsc_0_11_i_bcwt_drv;
  butterFly2_11_tw_h_butterFly2_11_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_11_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_11_i_s_raddr_core_sct);
  twiddle_h_rsc_0_11_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_11_tw_h_butterFly2_11_tw_h_and_nl));
  twiddle_h_rsc_0_11_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_11_i_s_din, twiddle_h_rsc_0_11_i_s_din_bfwt,
      twiddle_h_rsc_0_11_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_11_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_11_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_11_i_bcwt_drv OR
            twiddle_h_rsc_0_11_i_biwt)) OR twiddle_h_rsc_0_11_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_11_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_11_i_s_din_bfwt <= twiddle_h_rsc_0_11_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_11_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_11_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_11_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_11_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_11_i_bdwt <= twiddle_h_rsc_0_11_i_oswt AND core_wen;
  twiddle_h_rsc_0_11_i_biwt <= twiddle_h_rsc_0_11_i_ogwt AND twiddle_h_rsc_0_11_i_s_rrdy;
  twiddle_h_rsc_0_11_i_ogwt <= twiddle_h_rsc_0_11_i_oswt AND (NOT twiddle_h_rsc_0_11_i_bcwt);
  twiddle_h_rsc_0_11_i_s_re_core_sct <= twiddle_h_rsc_0_11_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_10_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_10_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_10_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_10_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_10_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_10_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_10_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_10_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp
    IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_10_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_10_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_10_tw_h_butterFly2_10_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_10_i_bcwt <= twiddle_h_rsc_0_10_i_bcwt_drv;

  twiddle_h_rsc_0_10_i_wen_comp <= (NOT twiddle_h_rsc_0_10_i_oswt) OR twiddle_h_rsc_0_10_i_biwt
      OR twiddle_h_rsc_0_10_i_bcwt_drv;
  butterFly2_10_tw_h_butterFly2_10_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_10_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_10_i_s_raddr_core_sct);
  twiddle_h_rsc_0_10_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_10_tw_h_butterFly2_10_tw_h_and_nl));
  twiddle_h_rsc_0_10_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_10_i_s_din, twiddle_h_rsc_0_10_i_s_din_bfwt,
      twiddle_h_rsc_0_10_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_10_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_10_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_10_i_bcwt_drv OR
            twiddle_h_rsc_0_10_i_biwt)) OR twiddle_h_rsc_0_10_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_10_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_10_i_s_din_bfwt <= twiddle_h_rsc_0_10_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_10_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_10_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_10_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_10_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_10_i_bdwt <= twiddle_h_rsc_0_10_i_oswt AND core_wen;
  twiddle_h_rsc_0_10_i_biwt <= twiddle_h_rsc_0_10_i_ogwt AND twiddle_h_rsc_0_10_i_s_rrdy;
  twiddle_h_rsc_0_10_i_ogwt <= twiddle_h_rsc_0_10_i_oswt AND (NOT twiddle_h_rsc_0_10_i_bcwt);
  twiddle_h_rsc_0_10_i_s_re_core_sct <= twiddle_h_rsc_0_10_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_9_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_9_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_9_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_9_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_9_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_9_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_9_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_9_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_9_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_9_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_9_tw_h_butterFly2_9_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_9_i_bcwt <= twiddle_h_rsc_0_9_i_bcwt_drv;

  twiddle_h_rsc_0_9_i_wen_comp <= (NOT twiddle_h_rsc_0_9_i_oswt) OR twiddle_h_rsc_0_9_i_biwt
      OR twiddle_h_rsc_0_9_i_bcwt_drv;
  butterFly2_9_tw_h_butterFly2_9_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_9_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_9_i_s_raddr_core_sct);
  twiddle_h_rsc_0_9_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_9_tw_h_butterFly2_9_tw_h_and_nl));
  twiddle_h_rsc_0_9_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_9_i_s_din, twiddle_h_rsc_0_9_i_s_din_bfwt,
      twiddle_h_rsc_0_9_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_9_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_9_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_9_i_bcwt_drv OR
            twiddle_h_rsc_0_9_i_biwt)) OR twiddle_h_rsc_0_9_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_9_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_9_i_s_din_bfwt <= twiddle_h_rsc_0_9_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_9_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_9_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_9_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_9_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_9_i_bdwt <= twiddle_h_rsc_0_9_i_oswt AND core_wen;
  twiddle_h_rsc_0_9_i_biwt <= twiddle_h_rsc_0_9_i_ogwt AND twiddle_h_rsc_0_9_i_s_rrdy;
  twiddle_h_rsc_0_9_i_ogwt <= twiddle_h_rsc_0_9_i_oswt AND (NOT twiddle_h_rsc_0_9_i_bcwt);
  twiddle_h_rsc_0_9_i_s_re_core_sct <= twiddle_h_rsc_0_9_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_8_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_8_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_8_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_8_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_8_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_8_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_8_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_8_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_8_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_8_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_8_tw_h_butterFly2_8_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_8_i_bcwt <= twiddle_h_rsc_0_8_i_bcwt_drv;

  twiddle_h_rsc_0_8_i_wen_comp <= (NOT twiddle_h_rsc_0_8_i_oswt) OR twiddle_h_rsc_0_8_i_biwt
      OR twiddle_h_rsc_0_8_i_bcwt_drv;
  butterFly2_8_tw_h_butterFly2_8_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_8_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_8_i_s_raddr_core_sct);
  twiddle_h_rsc_0_8_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_8_tw_h_butterFly2_8_tw_h_and_nl));
  twiddle_h_rsc_0_8_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_8_i_s_din, twiddle_h_rsc_0_8_i_s_din_bfwt,
      twiddle_h_rsc_0_8_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_8_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_8_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_8_i_bcwt_drv OR
            twiddle_h_rsc_0_8_i_biwt)) OR twiddle_h_rsc_0_8_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_8_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_8_i_s_din_bfwt <= twiddle_h_rsc_0_8_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_8_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_8_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_8_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_8_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_8_i_bdwt <= twiddle_h_rsc_0_8_i_oswt AND core_wen;
  twiddle_h_rsc_0_8_i_biwt <= twiddle_h_rsc_0_8_i_ogwt AND twiddle_h_rsc_0_8_i_s_rrdy;
  twiddle_h_rsc_0_8_i_ogwt <= twiddle_h_rsc_0_8_i_oswt AND (NOT twiddle_h_rsc_0_8_i_bcwt);
  twiddle_h_rsc_0_8_i_s_re_core_sct <= twiddle_h_rsc_0_8_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_7_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_7_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_7_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_7_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_7_tw_h_butterFly2_7_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_7_i_bcwt <= twiddle_h_rsc_0_7_i_bcwt_drv;

  twiddle_h_rsc_0_7_i_wen_comp <= (NOT twiddle_h_rsc_0_7_i_oswt) OR twiddle_h_rsc_0_7_i_biwt
      OR twiddle_h_rsc_0_7_i_bcwt_drv;
  butterFly2_7_tw_h_butterFly2_7_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_7_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_7_i_s_raddr_core_sct);
  twiddle_h_rsc_0_7_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_7_tw_h_butterFly2_7_tw_h_and_nl));
  twiddle_h_rsc_0_7_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_7_i_s_din, twiddle_h_rsc_0_7_i_s_din_bfwt,
      twiddle_h_rsc_0_7_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_7_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_7_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_7_i_bcwt_drv OR
            twiddle_h_rsc_0_7_i_biwt)) OR twiddle_h_rsc_0_7_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_7_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_7_i_s_din_bfwt <= twiddle_h_rsc_0_7_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_7_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_7_i_bdwt <= twiddle_h_rsc_0_7_i_oswt AND core_wen;
  twiddle_h_rsc_0_7_i_biwt <= twiddle_h_rsc_0_7_i_ogwt AND twiddle_h_rsc_0_7_i_s_rrdy;
  twiddle_h_rsc_0_7_i_ogwt <= twiddle_h_rsc_0_7_i_oswt AND (NOT twiddle_h_rsc_0_7_i_bcwt);
  twiddle_h_rsc_0_7_i_s_re_core_sct <= twiddle_h_rsc_0_7_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_6_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_6_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_6_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_6_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_6_tw_h_butterFly2_6_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_6_i_bcwt <= twiddle_h_rsc_0_6_i_bcwt_drv;

  twiddle_h_rsc_0_6_i_wen_comp <= (NOT twiddle_h_rsc_0_6_i_oswt) OR twiddle_h_rsc_0_6_i_biwt
      OR twiddle_h_rsc_0_6_i_bcwt_drv;
  butterFly2_6_tw_h_butterFly2_6_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_6_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_6_i_s_raddr_core_sct);
  twiddle_h_rsc_0_6_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_6_tw_h_butterFly2_6_tw_h_and_nl));
  twiddle_h_rsc_0_6_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_6_i_s_din, twiddle_h_rsc_0_6_i_s_din_bfwt,
      twiddle_h_rsc_0_6_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_6_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_6_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_6_i_bcwt_drv OR
            twiddle_h_rsc_0_6_i_biwt)) OR twiddle_h_rsc_0_6_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_6_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_6_i_s_din_bfwt <= twiddle_h_rsc_0_6_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_6_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_6_i_bdwt <= twiddle_h_rsc_0_6_i_oswt AND core_wen;
  twiddle_h_rsc_0_6_i_biwt <= twiddle_h_rsc_0_6_i_ogwt AND twiddle_h_rsc_0_6_i_s_rrdy;
  twiddle_h_rsc_0_6_i_ogwt <= twiddle_h_rsc_0_6_i_oswt AND (NOT twiddle_h_rsc_0_6_i_bcwt);
  twiddle_h_rsc_0_6_i_s_re_core_sct <= twiddle_h_rsc_0_6_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_5_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_5_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_5_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_5_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_5_tw_h_butterFly2_5_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_5_i_bcwt <= twiddle_h_rsc_0_5_i_bcwt_drv;

  twiddle_h_rsc_0_5_i_wen_comp <= (NOT twiddle_h_rsc_0_5_i_oswt) OR twiddle_h_rsc_0_5_i_biwt
      OR twiddle_h_rsc_0_5_i_bcwt_drv;
  butterFly2_5_tw_h_butterFly2_5_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_5_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_5_i_s_raddr_core_sct);
  twiddle_h_rsc_0_5_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_5_tw_h_butterFly2_5_tw_h_and_nl));
  twiddle_h_rsc_0_5_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_5_i_s_din, twiddle_h_rsc_0_5_i_s_din_bfwt,
      twiddle_h_rsc_0_5_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_5_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_5_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_5_i_bcwt_drv OR
            twiddle_h_rsc_0_5_i_biwt)) OR twiddle_h_rsc_0_5_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_5_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_5_i_s_din_bfwt <= twiddle_h_rsc_0_5_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_5_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_5_i_bdwt <= twiddle_h_rsc_0_5_i_oswt AND core_wen;
  twiddle_h_rsc_0_5_i_biwt <= twiddle_h_rsc_0_5_i_ogwt AND twiddle_h_rsc_0_5_i_s_rrdy;
  twiddle_h_rsc_0_5_i_ogwt <= twiddle_h_rsc_0_5_i_oswt AND (NOT twiddle_h_rsc_0_5_i_bcwt);
  twiddle_h_rsc_0_5_i_s_re_core_sct <= twiddle_h_rsc_0_5_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_4_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_4_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_4_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_4_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_4_tw_h_butterFly2_4_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_4_i_bcwt <= twiddle_h_rsc_0_4_i_bcwt_drv;

  twiddle_h_rsc_0_4_i_wen_comp <= (NOT twiddle_h_rsc_0_4_i_oswt) OR twiddle_h_rsc_0_4_i_biwt
      OR twiddle_h_rsc_0_4_i_bcwt_drv;
  butterFly2_4_tw_h_butterFly2_4_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_4_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_4_i_s_raddr_core_sct);
  twiddle_h_rsc_0_4_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_4_tw_h_butterFly2_4_tw_h_and_nl));
  twiddle_h_rsc_0_4_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_4_i_s_din, twiddle_h_rsc_0_4_i_s_din_bfwt,
      twiddle_h_rsc_0_4_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_4_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_4_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_4_i_bcwt_drv OR
            twiddle_h_rsc_0_4_i_biwt)) OR twiddle_h_rsc_0_4_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_4_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_4_i_s_din_bfwt <= twiddle_h_rsc_0_4_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_4_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_4_i_bdwt <= twiddle_h_rsc_0_4_i_oswt AND core_wen;
  twiddle_h_rsc_0_4_i_biwt <= twiddle_h_rsc_0_4_i_ogwt AND twiddle_h_rsc_0_4_i_s_rrdy;
  twiddle_h_rsc_0_4_i_ogwt <= twiddle_h_rsc_0_4_i_oswt AND (NOT twiddle_h_rsc_0_4_i_bcwt);
  twiddle_h_rsc_0_4_i_s_re_core_sct <= twiddle_h_rsc_0_4_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_3_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_3_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_3_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_3_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_3_tw_h_butterFly2_3_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_3_i_bcwt <= twiddle_h_rsc_0_3_i_bcwt_drv;

  twiddle_h_rsc_0_3_i_wen_comp <= (NOT twiddle_h_rsc_0_3_i_oswt) OR twiddle_h_rsc_0_3_i_biwt
      OR twiddle_h_rsc_0_3_i_bcwt_drv;
  butterFly2_3_tw_h_butterFly2_3_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_3_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_3_i_s_raddr_core_sct);
  twiddle_h_rsc_0_3_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_3_tw_h_butterFly2_3_tw_h_and_nl));
  twiddle_h_rsc_0_3_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_3_i_s_din, twiddle_h_rsc_0_3_i_s_din_bfwt,
      twiddle_h_rsc_0_3_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_3_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_3_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_3_i_bcwt_drv OR
            twiddle_h_rsc_0_3_i_biwt)) OR twiddle_h_rsc_0_3_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_3_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_3_i_s_din_bfwt <= twiddle_h_rsc_0_3_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_3_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_3_i_bdwt <= twiddle_h_rsc_0_3_i_oswt AND core_wen;
  twiddle_h_rsc_0_3_i_biwt <= twiddle_h_rsc_0_3_i_ogwt AND twiddle_h_rsc_0_3_i_s_rrdy;
  twiddle_h_rsc_0_3_i_ogwt <= twiddle_h_rsc_0_3_i_oswt AND (NOT twiddle_h_rsc_0_3_i_bcwt);
  twiddle_h_rsc_0_3_i_s_re_core_sct <= twiddle_h_rsc_0_3_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_2_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_2_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_2_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_2_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_2_tw_h_butterFly2_2_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_2_i_bcwt <= twiddle_h_rsc_0_2_i_bcwt_drv;

  twiddle_h_rsc_0_2_i_wen_comp <= (NOT twiddle_h_rsc_0_2_i_oswt) OR twiddle_h_rsc_0_2_i_biwt
      OR twiddle_h_rsc_0_2_i_bcwt_drv;
  butterFly2_2_tw_h_butterFly2_2_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_2_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_2_i_s_raddr_core_sct);
  twiddle_h_rsc_0_2_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_2_tw_h_butterFly2_2_tw_h_and_nl));
  twiddle_h_rsc_0_2_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_2_i_s_din, twiddle_h_rsc_0_2_i_s_din_bfwt,
      twiddle_h_rsc_0_2_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_2_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_2_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_2_i_bcwt_drv OR
            twiddle_h_rsc_0_2_i_biwt)) OR twiddle_h_rsc_0_2_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_2_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_2_i_s_din_bfwt <= twiddle_h_rsc_0_2_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_2_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_2_i_bdwt <= twiddle_h_rsc_0_2_i_oswt AND core_wen;
  twiddle_h_rsc_0_2_i_biwt <= twiddle_h_rsc_0_2_i_ogwt AND twiddle_h_rsc_0_2_i_s_rrdy;
  twiddle_h_rsc_0_2_i_ogwt <= twiddle_h_rsc_0_2_i_oswt AND (NOT twiddle_h_rsc_0_2_i_bcwt);
  twiddle_h_rsc_0_2_i_s_re_core_sct <= twiddle_h_rsc_0_2_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_1_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_1_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_1_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_1_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_1_tw_h_butterFly2_1_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_1_i_bcwt <= twiddle_h_rsc_0_1_i_bcwt_drv;

  twiddle_h_rsc_0_1_i_wen_comp <= (NOT twiddle_h_rsc_0_1_i_oswt) OR twiddle_h_rsc_0_1_i_biwt
      OR twiddle_h_rsc_0_1_i_bcwt_drv;
  butterFly2_1_tw_h_butterFly2_1_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_1_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_1_i_s_raddr_core_sct);
  twiddle_h_rsc_0_1_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_1_tw_h_butterFly2_1_tw_h_and_nl));
  twiddle_h_rsc_0_1_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_1_i_s_din, twiddle_h_rsc_0_1_i_s_din_bfwt,
      twiddle_h_rsc_0_1_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_1_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_1_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_1_i_bcwt_drv OR
            twiddle_h_rsc_0_1_i_biwt)) OR twiddle_h_rsc_0_1_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_1_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_1_i_s_din_bfwt <= twiddle_h_rsc_0_1_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_1_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_1_i_bdwt <= twiddle_h_rsc_0_1_i_oswt AND core_wen;
  twiddle_h_rsc_0_1_i_biwt <= twiddle_h_rsc_0_1_i_ogwt AND twiddle_h_rsc_0_1_i_s_rrdy;
  twiddle_h_rsc_0_1_i_ogwt <= twiddle_h_rsc_0_1_i_oswt AND (NOT twiddle_h_rsc_0_1_i_bcwt);
  twiddle_h_rsc_0_1_i_s_re_core_sct <= twiddle_h_rsc_0_1_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_i_biwt : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_bdwt : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_bcwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_0_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_h_rsc_0_0_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL INNER_LOOP1_tw_h_INNER_LOOP1_tw_h_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_h_rsc_0_0_i_bcwt <= twiddle_h_rsc_0_0_i_bcwt_drv;

  twiddle_h_rsc_0_0_i_wen_comp <= (NOT twiddle_h_rsc_0_0_i_oswt) OR twiddle_h_rsc_0_0_i_biwt
      OR twiddle_h_rsc_0_0_i_bcwt_drv;
  INNER_LOOP1_tw_h_INNER_LOOP1_tw_h_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_h_rsc_0_0_i_s_raddr_core(4 DOWNTO 0)), twiddle_h_rsc_0_0_i_s_raddr_core_sct);
  twiddle_h_rsc_0_0_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(INNER_LOOP1_tw_h_INNER_LOOP1_tw_h_and_nl));
  twiddle_h_rsc_0_0_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_h_rsc_0_0_i_s_din, twiddle_h_rsc_0_0_i_s_din_bfwt,
      twiddle_h_rsc_0_0_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_h_rsc_0_0_i_bcwt_drv <= '0';
      ELSE
        twiddle_h_rsc_0_0_i_bcwt_drv <= NOT((NOT(twiddle_h_rsc_0_0_i_bcwt_drv OR
            twiddle_h_rsc_0_0_i_biwt)) OR twiddle_h_rsc_0_0_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_h_rsc_0_0_i_biwt = '1' ) THEN
        twiddle_h_rsc_0_0_i_s_din_bfwt <= twiddle_h_rsc_0_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_biwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_i_bdwt : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_i_bcwt : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_ctrl
    IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_0_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_h_rsc_0_0_i_bdwt <= twiddle_h_rsc_0_0_i_oswt AND core_wen;
  twiddle_h_rsc_0_0_i_biwt <= twiddle_h_rsc_0_0_i_ogwt AND twiddle_h_rsc_0_0_i_s_rrdy;
  twiddle_h_rsc_0_0_i_ogwt <= twiddle_h_rsc_0_0_i_oswt AND (NOT twiddle_h_rsc_0_0_i_bcwt);
  twiddle_h_rsc_0_0_i_s_re_core_sct <= twiddle_h_rsc_0_0_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_15_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_15_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_15_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_15_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_15_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_15_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_15_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_15_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_15_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_15_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_15_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_15_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_15_tw_butterFly2_15_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_15_i_bcwt <= twiddle_rsc_0_15_i_bcwt_drv;

  twiddle_rsc_0_15_i_wen_comp <= (NOT twiddle_rsc_0_15_i_oswt) OR twiddle_rsc_0_15_i_biwt
      OR twiddle_rsc_0_15_i_bcwt_drv;
  butterFly2_15_tw_butterFly2_15_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_15_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_15_i_s_raddr_core_sct);
  twiddle_rsc_0_15_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_15_tw_butterFly2_15_tw_and_nl));
  twiddle_rsc_0_15_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_15_i_s_din, twiddle_rsc_0_15_i_s_din_bfwt,
      twiddle_rsc_0_15_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_15_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_15_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_15_i_bcwt_drv OR twiddle_rsc_0_15_i_biwt))
            OR twiddle_rsc_0_15_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_15_i_biwt = '1' ) THEN
        twiddle_rsc_0_15_i_s_din_bfwt <= twiddle_rsc_0_15_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_15_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_15_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_15_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_15_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_15_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_15_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_15_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_15_i_bdwt <= twiddle_rsc_0_15_i_oswt AND core_wen;
  twiddle_rsc_0_15_i_biwt <= twiddle_rsc_0_15_i_ogwt AND twiddle_rsc_0_15_i_s_rrdy;
  twiddle_rsc_0_15_i_ogwt <= twiddle_rsc_0_15_i_oswt AND (NOT twiddle_rsc_0_15_i_bcwt);
  twiddle_rsc_0_15_i_s_re_core_sct <= twiddle_rsc_0_15_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_14_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_14_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_14_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_14_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_14_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_14_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_14_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_14_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_14_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_14_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_14_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_14_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_14_tw_butterFly2_14_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_14_i_bcwt <= twiddle_rsc_0_14_i_bcwt_drv;

  twiddle_rsc_0_14_i_wen_comp <= (NOT twiddle_rsc_0_14_i_oswt) OR twiddle_rsc_0_14_i_biwt
      OR twiddle_rsc_0_14_i_bcwt_drv;
  butterFly2_14_tw_butterFly2_14_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_14_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_14_i_s_raddr_core_sct);
  twiddle_rsc_0_14_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_14_tw_butterFly2_14_tw_and_nl));
  twiddle_rsc_0_14_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_14_i_s_din, twiddle_rsc_0_14_i_s_din_bfwt,
      twiddle_rsc_0_14_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_14_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_14_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_14_i_bcwt_drv OR twiddle_rsc_0_14_i_biwt))
            OR twiddle_rsc_0_14_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_14_i_biwt = '1' ) THEN
        twiddle_rsc_0_14_i_s_din_bfwt <= twiddle_rsc_0_14_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_14_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_14_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_14_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_14_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_14_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_14_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_14_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_14_i_bdwt <= twiddle_rsc_0_14_i_oswt AND core_wen;
  twiddle_rsc_0_14_i_biwt <= twiddle_rsc_0_14_i_ogwt AND twiddle_rsc_0_14_i_s_rrdy;
  twiddle_rsc_0_14_i_ogwt <= twiddle_rsc_0_14_i_oswt AND (NOT twiddle_rsc_0_14_i_bcwt);
  twiddle_rsc_0_14_i_s_re_core_sct <= twiddle_rsc_0_14_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_13_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_13_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_13_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_13_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_13_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_13_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_13_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_13_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_13_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_13_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_13_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_13_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_13_tw_butterFly2_13_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_13_i_bcwt <= twiddle_rsc_0_13_i_bcwt_drv;

  twiddle_rsc_0_13_i_wen_comp <= (NOT twiddle_rsc_0_13_i_oswt) OR twiddle_rsc_0_13_i_biwt
      OR twiddle_rsc_0_13_i_bcwt_drv;
  butterFly2_13_tw_butterFly2_13_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_13_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_13_i_s_raddr_core_sct);
  twiddle_rsc_0_13_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_13_tw_butterFly2_13_tw_and_nl));
  twiddle_rsc_0_13_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_13_i_s_din, twiddle_rsc_0_13_i_s_din_bfwt,
      twiddle_rsc_0_13_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_13_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_13_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_13_i_bcwt_drv OR twiddle_rsc_0_13_i_biwt))
            OR twiddle_rsc_0_13_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_13_i_biwt = '1' ) THEN
        twiddle_rsc_0_13_i_s_din_bfwt <= twiddle_rsc_0_13_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_13_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_13_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_13_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_13_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_13_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_13_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_13_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_13_i_bdwt <= twiddle_rsc_0_13_i_oswt AND core_wen;
  twiddle_rsc_0_13_i_biwt <= twiddle_rsc_0_13_i_ogwt AND twiddle_rsc_0_13_i_s_rrdy;
  twiddle_rsc_0_13_i_ogwt <= twiddle_rsc_0_13_i_oswt AND (NOT twiddle_rsc_0_13_i_bcwt);
  twiddle_rsc_0_13_i_s_re_core_sct <= twiddle_rsc_0_13_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_12_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_12_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_12_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_12_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_12_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_12_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_12_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_12_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_12_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_12_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_12_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_12_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_12_tw_butterFly2_12_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_12_i_bcwt <= twiddle_rsc_0_12_i_bcwt_drv;

  twiddle_rsc_0_12_i_wen_comp <= (NOT twiddle_rsc_0_12_i_oswt) OR twiddle_rsc_0_12_i_biwt
      OR twiddle_rsc_0_12_i_bcwt_drv;
  butterFly2_12_tw_butterFly2_12_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_12_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_12_i_s_raddr_core_sct);
  twiddle_rsc_0_12_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_12_tw_butterFly2_12_tw_and_nl));
  twiddle_rsc_0_12_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_12_i_s_din, twiddle_rsc_0_12_i_s_din_bfwt,
      twiddle_rsc_0_12_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_12_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_12_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_12_i_bcwt_drv OR twiddle_rsc_0_12_i_biwt))
            OR twiddle_rsc_0_12_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_12_i_biwt = '1' ) THEN
        twiddle_rsc_0_12_i_s_din_bfwt <= twiddle_rsc_0_12_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_12_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_12_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_12_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_12_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_12_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_12_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_12_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_12_i_bdwt <= twiddle_rsc_0_12_i_oswt AND core_wen;
  twiddle_rsc_0_12_i_biwt <= twiddle_rsc_0_12_i_ogwt AND twiddle_rsc_0_12_i_s_rrdy;
  twiddle_rsc_0_12_i_ogwt <= twiddle_rsc_0_12_i_oswt AND (NOT twiddle_rsc_0_12_i_bcwt);
  twiddle_rsc_0_12_i_s_re_core_sct <= twiddle_rsc_0_12_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_11_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_11_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_11_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_11_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_11_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_11_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_11_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_11_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_11_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_11_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_11_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_11_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_11_tw_butterFly2_11_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_11_i_bcwt <= twiddle_rsc_0_11_i_bcwt_drv;

  twiddle_rsc_0_11_i_wen_comp <= (NOT twiddle_rsc_0_11_i_oswt) OR twiddle_rsc_0_11_i_biwt
      OR twiddle_rsc_0_11_i_bcwt_drv;
  butterFly2_11_tw_butterFly2_11_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_11_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_11_i_s_raddr_core_sct);
  twiddle_rsc_0_11_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_11_tw_butterFly2_11_tw_and_nl));
  twiddle_rsc_0_11_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_11_i_s_din, twiddle_rsc_0_11_i_s_din_bfwt,
      twiddle_rsc_0_11_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_11_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_11_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_11_i_bcwt_drv OR twiddle_rsc_0_11_i_biwt))
            OR twiddle_rsc_0_11_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_11_i_biwt = '1' ) THEN
        twiddle_rsc_0_11_i_s_din_bfwt <= twiddle_rsc_0_11_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_11_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_11_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_11_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_11_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_11_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_11_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_11_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_11_i_bdwt <= twiddle_rsc_0_11_i_oswt AND core_wen;
  twiddle_rsc_0_11_i_biwt <= twiddle_rsc_0_11_i_ogwt AND twiddle_rsc_0_11_i_s_rrdy;
  twiddle_rsc_0_11_i_ogwt <= twiddle_rsc_0_11_i_oswt AND (NOT twiddle_rsc_0_11_i_bcwt);
  twiddle_rsc_0_11_i_s_re_core_sct <= twiddle_rsc_0_11_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_10_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_10_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_10_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_10_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_10_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_10_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_10_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_10_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_10_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_10_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_10_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_10_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_10_tw_butterFly2_10_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_10_i_bcwt <= twiddle_rsc_0_10_i_bcwt_drv;

  twiddle_rsc_0_10_i_wen_comp <= (NOT twiddle_rsc_0_10_i_oswt) OR twiddle_rsc_0_10_i_biwt
      OR twiddle_rsc_0_10_i_bcwt_drv;
  butterFly2_10_tw_butterFly2_10_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_10_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_10_i_s_raddr_core_sct);
  twiddle_rsc_0_10_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_10_tw_butterFly2_10_tw_and_nl));
  twiddle_rsc_0_10_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_10_i_s_din, twiddle_rsc_0_10_i_s_din_bfwt,
      twiddle_rsc_0_10_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_10_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_10_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_10_i_bcwt_drv OR twiddle_rsc_0_10_i_biwt))
            OR twiddle_rsc_0_10_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_10_i_biwt = '1' ) THEN
        twiddle_rsc_0_10_i_s_din_bfwt <= twiddle_rsc_0_10_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_10_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_10_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_10_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_10_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_10_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_10_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_10_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_10_i_bdwt <= twiddle_rsc_0_10_i_oswt AND core_wen;
  twiddle_rsc_0_10_i_biwt <= twiddle_rsc_0_10_i_ogwt AND twiddle_rsc_0_10_i_s_rrdy;
  twiddle_rsc_0_10_i_ogwt <= twiddle_rsc_0_10_i_oswt AND (NOT twiddle_rsc_0_10_i_bcwt);
  twiddle_rsc_0_10_i_s_re_core_sct <= twiddle_rsc_0_10_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_9_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_9_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_9_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_9_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_9_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_9_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_9_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_9_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_9_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_9_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_9_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_9_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_9_tw_butterFly2_9_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_9_i_bcwt <= twiddle_rsc_0_9_i_bcwt_drv;

  twiddle_rsc_0_9_i_wen_comp <= (NOT twiddle_rsc_0_9_i_oswt) OR twiddle_rsc_0_9_i_biwt
      OR twiddle_rsc_0_9_i_bcwt_drv;
  butterFly2_9_tw_butterFly2_9_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_9_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_9_i_s_raddr_core_sct);
  twiddle_rsc_0_9_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_9_tw_butterFly2_9_tw_and_nl));
  twiddle_rsc_0_9_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_9_i_s_din, twiddle_rsc_0_9_i_s_din_bfwt,
      twiddle_rsc_0_9_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_9_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_9_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_9_i_bcwt_drv OR twiddle_rsc_0_9_i_biwt))
            OR twiddle_rsc_0_9_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_9_i_biwt = '1' ) THEN
        twiddle_rsc_0_9_i_s_din_bfwt <= twiddle_rsc_0_9_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_9_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_9_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_9_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_9_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_9_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_9_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_9_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_9_i_bdwt <= twiddle_rsc_0_9_i_oswt AND core_wen;
  twiddle_rsc_0_9_i_biwt <= twiddle_rsc_0_9_i_ogwt AND twiddle_rsc_0_9_i_s_rrdy;
  twiddle_rsc_0_9_i_ogwt <= twiddle_rsc_0_9_i_oswt AND (NOT twiddle_rsc_0_9_i_bcwt);
  twiddle_rsc_0_9_i_s_re_core_sct <= twiddle_rsc_0_9_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_8_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_8_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_8_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_8_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_8_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_8_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_8_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_8_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_8_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_8_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_8_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_8_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_8_tw_butterFly2_8_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_8_i_bcwt <= twiddle_rsc_0_8_i_bcwt_drv;

  twiddle_rsc_0_8_i_wen_comp <= (NOT twiddle_rsc_0_8_i_oswt) OR twiddle_rsc_0_8_i_biwt
      OR twiddle_rsc_0_8_i_bcwt_drv;
  butterFly2_8_tw_butterFly2_8_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_8_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_8_i_s_raddr_core_sct);
  twiddle_rsc_0_8_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_8_tw_butterFly2_8_tw_and_nl));
  twiddle_rsc_0_8_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_8_i_s_din, twiddle_rsc_0_8_i_s_din_bfwt,
      twiddle_rsc_0_8_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_8_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_8_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_8_i_bcwt_drv OR twiddle_rsc_0_8_i_biwt))
            OR twiddle_rsc_0_8_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_8_i_biwt = '1' ) THEN
        twiddle_rsc_0_8_i_s_din_bfwt <= twiddle_rsc_0_8_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_8_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_8_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_8_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_8_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_8_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_8_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_8_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_8_i_bdwt <= twiddle_rsc_0_8_i_oswt AND core_wen;
  twiddle_rsc_0_8_i_biwt <= twiddle_rsc_0_8_i_ogwt AND twiddle_rsc_0_8_i_s_rrdy;
  twiddle_rsc_0_8_i_ogwt <= twiddle_rsc_0_8_i_oswt AND (NOT twiddle_rsc_0_8_i_bcwt);
  twiddle_rsc_0_8_i_s_re_core_sct <= twiddle_rsc_0_8_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_7_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_7_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_7_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_7_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_7_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_7_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_7_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_7_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_7_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_7_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_7_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_7_tw_butterFly2_7_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_7_i_bcwt <= twiddle_rsc_0_7_i_bcwt_drv;

  twiddle_rsc_0_7_i_wen_comp <= (NOT twiddle_rsc_0_7_i_oswt) OR twiddle_rsc_0_7_i_biwt
      OR twiddle_rsc_0_7_i_bcwt_drv;
  butterFly2_7_tw_butterFly2_7_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_7_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_7_i_s_raddr_core_sct);
  twiddle_rsc_0_7_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_7_tw_butterFly2_7_tw_and_nl));
  twiddle_rsc_0_7_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_7_i_s_din, twiddle_rsc_0_7_i_s_din_bfwt,
      twiddle_rsc_0_7_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_7_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_7_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_7_i_bcwt_drv OR twiddle_rsc_0_7_i_biwt))
            OR twiddle_rsc_0_7_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_7_i_biwt = '1' ) THEN
        twiddle_rsc_0_7_i_s_din_bfwt <= twiddle_rsc_0_7_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_7_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_7_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_7_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_7_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_7_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_7_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_7_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_7_i_bdwt <= twiddle_rsc_0_7_i_oswt AND core_wen;
  twiddle_rsc_0_7_i_biwt <= twiddle_rsc_0_7_i_ogwt AND twiddle_rsc_0_7_i_s_rrdy;
  twiddle_rsc_0_7_i_ogwt <= twiddle_rsc_0_7_i_oswt AND (NOT twiddle_rsc_0_7_i_bcwt);
  twiddle_rsc_0_7_i_s_re_core_sct <= twiddle_rsc_0_7_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_6_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_6_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_6_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_6_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_6_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_6_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_6_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_6_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_6_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_6_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_6_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_6_tw_butterFly2_6_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_6_i_bcwt <= twiddle_rsc_0_6_i_bcwt_drv;

  twiddle_rsc_0_6_i_wen_comp <= (NOT twiddle_rsc_0_6_i_oswt) OR twiddle_rsc_0_6_i_biwt
      OR twiddle_rsc_0_6_i_bcwt_drv;
  butterFly2_6_tw_butterFly2_6_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_6_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_6_i_s_raddr_core_sct);
  twiddle_rsc_0_6_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_6_tw_butterFly2_6_tw_and_nl));
  twiddle_rsc_0_6_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_6_i_s_din, twiddle_rsc_0_6_i_s_din_bfwt,
      twiddle_rsc_0_6_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_6_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_6_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_6_i_bcwt_drv OR twiddle_rsc_0_6_i_biwt))
            OR twiddle_rsc_0_6_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_6_i_biwt = '1' ) THEN
        twiddle_rsc_0_6_i_s_din_bfwt <= twiddle_rsc_0_6_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_6_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_6_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_6_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_6_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_6_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_6_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_6_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_6_i_bdwt <= twiddle_rsc_0_6_i_oswt AND core_wen;
  twiddle_rsc_0_6_i_biwt <= twiddle_rsc_0_6_i_ogwt AND twiddle_rsc_0_6_i_s_rrdy;
  twiddle_rsc_0_6_i_ogwt <= twiddle_rsc_0_6_i_oswt AND (NOT twiddle_rsc_0_6_i_bcwt);
  twiddle_rsc_0_6_i_s_re_core_sct <= twiddle_rsc_0_6_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_5_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_5_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_5_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_5_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_5_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_5_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_5_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_5_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_5_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_5_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_5_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_5_tw_butterFly2_5_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_5_i_bcwt <= twiddle_rsc_0_5_i_bcwt_drv;

  twiddle_rsc_0_5_i_wen_comp <= (NOT twiddle_rsc_0_5_i_oswt) OR twiddle_rsc_0_5_i_biwt
      OR twiddle_rsc_0_5_i_bcwt_drv;
  butterFly2_5_tw_butterFly2_5_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_5_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_5_i_s_raddr_core_sct);
  twiddle_rsc_0_5_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_5_tw_butterFly2_5_tw_and_nl));
  twiddle_rsc_0_5_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_5_i_s_din, twiddle_rsc_0_5_i_s_din_bfwt,
      twiddle_rsc_0_5_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_5_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_5_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_5_i_bcwt_drv OR twiddle_rsc_0_5_i_biwt))
            OR twiddle_rsc_0_5_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_5_i_biwt = '1' ) THEN
        twiddle_rsc_0_5_i_s_din_bfwt <= twiddle_rsc_0_5_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_5_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_5_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_5_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_5_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_5_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_5_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_5_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_5_i_bdwt <= twiddle_rsc_0_5_i_oswt AND core_wen;
  twiddle_rsc_0_5_i_biwt <= twiddle_rsc_0_5_i_ogwt AND twiddle_rsc_0_5_i_s_rrdy;
  twiddle_rsc_0_5_i_ogwt <= twiddle_rsc_0_5_i_oswt AND (NOT twiddle_rsc_0_5_i_bcwt);
  twiddle_rsc_0_5_i_s_re_core_sct <= twiddle_rsc_0_5_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_4_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_4_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_4_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_4_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_4_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_4_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_4_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_4_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_4_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_4_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_4_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_4_tw_butterFly2_4_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_4_i_bcwt <= twiddle_rsc_0_4_i_bcwt_drv;

  twiddle_rsc_0_4_i_wen_comp <= (NOT twiddle_rsc_0_4_i_oswt) OR twiddle_rsc_0_4_i_biwt
      OR twiddle_rsc_0_4_i_bcwt_drv;
  butterFly2_4_tw_butterFly2_4_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_4_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_4_i_s_raddr_core_sct);
  twiddle_rsc_0_4_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_4_tw_butterFly2_4_tw_and_nl));
  twiddle_rsc_0_4_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_4_i_s_din, twiddle_rsc_0_4_i_s_din_bfwt,
      twiddle_rsc_0_4_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_4_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_4_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_4_i_bcwt_drv OR twiddle_rsc_0_4_i_biwt))
            OR twiddle_rsc_0_4_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_4_i_biwt = '1' ) THEN
        twiddle_rsc_0_4_i_s_din_bfwt <= twiddle_rsc_0_4_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_4_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_4_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_4_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_4_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_4_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_4_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_4_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_4_i_bdwt <= twiddle_rsc_0_4_i_oswt AND core_wen;
  twiddle_rsc_0_4_i_biwt <= twiddle_rsc_0_4_i_ogwt AND twiddle_rsc_0_4_i_s_rrdy;
  twiddle_rsc_0_4_i_ogwt <= twiddle_rsc_0_4_i_oswt AND (NOT twiddle_rsc_0_4_i_bcwt);
  twiddle_rsc_0_4_i_s_re_core_sct <= twiddle_rsc_0_4_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_3_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_3_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_3_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_3_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_3_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_3_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_3_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_3_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_3_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_3_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_3_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_3_tw_butterFly2_3_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_3_i_bcwt <= twiddle_rsc_0_3_i_bcwt_drv;

  twiddle_rsc_0_3_i_wen_comp <= (NOT twiddle_rsc_0_3_i_oswt) OR twiddle_rsc_0_3_i_biwt
      OR twiddle_rsc_0_3_i_bcwt_drv;
  butterFly2_3_tw_butterFly2_3_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_3_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_3_i_s_raddr_core_sct);
  twiddle_rsc_0_3_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_3_tw_butterFly2_3_tw_and_nl));
  twiddle_rsc_0_3_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_3_i_s_din, twiddle_rsc_0_3_i_s_din_bfwt,
      twiddle_rsc_0_3_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_3_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_3_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_3_i_bcwt_drv OR twiddle_rsc_0_3_i_biwt))
            OR twiddle_rsc_0_3_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_3_i_biwt = '1' ) THEN
        twiddle_rsc_0_3_i_s_din_bfwt <= twiddle_rsc_0_3_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_3_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_3_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_3_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_3_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_3_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_3_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_3_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_3_i_bdwt <= twiddle_rsc_0_3_i_oswt AND core_wen;
  twiddle_rsc_0_3_i_biwt <= twiddle_rsc_0_3_i_ogwt AND twiddle_rsc_0_3_i_s_rrdy;
  twiddle_rsc_0_3_i_ogwt <= twiddle_rsc_0_3_i_oswt AND (NOT twiddle_rsc_0_3_i_bcwt);
  twiddle_rsc_0_3_i_s_re_core_sct <= twiddle_rsc_0_3_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_2_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_2_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_2_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_2_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_2_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_2_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_2_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_2_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_2_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_2_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_2_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_2_tw_butterFly2_2_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_2_i_bcwt <= twiddle_rsc_0_2_i_bcwt_drv;

  twiddle_rsc_0_2_i_wen_comp <= (NOT twiddle_rsc_0_2_i_oswt) OR twiddle_rsc_0_2_i_biwt
      OR twiddle_rsc_0_2_i_bcwt_drv;
  butterFly2_2_tw_butterFly2_2_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_2_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_2_i_s_raddr_core_sct);
  twiddle_rsc_0_2_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_2_tw_butterFly2_2_tw_and_nl));
  twiddle_rsc_0_2_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_2_i_s_din, twiddle_rsc_0_2_i_s_din_bfwt,
      twiddle_rsc_0_2_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_2_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_2_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_2_i_bcwt_drv OR twiddle_rsc_0_2_i_biwt))
            OR twiddle_rsc_0_2_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_2_i_biwt = '1' ) THEN
        twiddle_rsc_0_2_i_s_din_bfwt <= twiddle_rsc_0_2_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_2_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_2_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_2_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_2_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_2_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_2_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_2_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_2_i_bdwt <= twiddle_rsc_0_2_i_oswt AND core_wen;
  twiddle_rsc_0_2_i_biwt <= twiddle_rsc_0_2_i_ogwt AND twiddle_rsc_0_2_i_s_rrdy;
  twiddle_rsc_0_2_i_ogwt <= twiddle_rsc_0_2_i_oswt AND (NOT twiddle_rsc_0_2_i_bcwt);
  twiddle_rsc_0_2_i_s_re_core_sct <= twiddle_rsc_0_2_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_1_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_1_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_1_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_1_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_1_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_1_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_1_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_1_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_1_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_1_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_1_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL butterFly2_1_tw_butterFly2_1_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_1_i_bcwt <= twiddle_rsc_0_1_i_bcwt_drv;

  twiddle_rsc_0_1_i_wen_comp <= (NOT twiddle_rsc_0_1_i_oswt) OR twiddle_rsc_0_1_i_biwt
      OR twiddle_rsc_0_1_i_bcwt_drv;
  butterFly2_1_tw_butterFly2_1_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_1_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_1_i_s_raddr_core_sct);
  twiddle_rsc_0_1_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(butterFly2_1_tw_butterFly2_1_tw_and_nl));
  twiddle_rsc_0_1_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_1_i_s_din, twiddle_rsc_0_1_i_s_din_bfwt,
      twiddle_rsc_0_1_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_1_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_1_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_1_i_bcwt_drv OR twiddle_rsc_0_1_i_biwt))
            OR twiddle_rsc_0_1_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_1_i_biwt = '1' ) THEN
        twiddle_rsc_0_1_i_s_din_bfwt <= twiddle_rsc_0_1_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_1_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_1_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_1_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_1_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_1_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_1_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_1_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_1_i_bdwt <= twiddle_rsc_0_1_i_oswt AND core_wen;
  twiddle_rsc_0_1_i_biwt <= twiddle_rsc_0_1_i_ogwt AND twiddle_rsc_0_1_i_s_rrdy;
  twiddle_rsc_0_1_i_ogwt <= twiddle_rsc_0_1_i_oswt AND (NOT twiddle_rsc_0_1_i_bcwt);
  twiddle_rsc_0_1_i_s_re_core_sct <= twiddle_rsc_0_1_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_0_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_0_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_i_biwt : IN STD_LOGIC;
    twiddle_rsc_0_0_i_bdwt : IN STD_LOGIC;
    twiddle_rsc_0_0_i_bcwt : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_0_i_s_raddr_core_sct : IN STD_LOGIC;
    twiddle_rsc_0_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp IS
  -- Default Constants

  -- Output Reader Declarations
  SIGNAL twiddle_rsc_0_0_i_bcwt_drv : STD_LOGIC;

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_0_i_s_din_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL INNER_LOOP1_tw_INNER_LOOP1_tw_and_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  -- Output Reader Assignments
  twiddle_rsc_0_0_i_bcwt <= twiddle_rsc_0_0_i_bcwt_drv;

  twiddle_rsc_0_0_i_wen_comp <= (NOT twiddle_rsc_0_0_i_oswt) OR twiddle_rsc_0_0_i_biwt
      OR twiddle_rsc_0_0_i_bcwt_drv;
  INNER_LOOP1_tw_INNER_LOOP1_tw_and_nl <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (twiddle_rsc_0_0_i_s_raddr_core(4 DOWNTO 0)), twiddle_rsc_0_0_i_s_raddr_core_sct);
  twiddle_rsc_0_0_i_s_raddr <= STD_LOGIC_VECTOR(UNSIGNED'( "0") & UNSIGNED(INNER_LOOP1_tw_INNER_LOOP1_tw_and_nl));
  twiddle_rsc_0_0_i_s_din_mxwt <= MUX_v_32_2_2(twiddle_rsc_0_0_i_s_din, twiddle_rsc_0_0_i_s_din_bfwt,
      twiddle_rsc_0_0_i_bcwt_drv);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        twiddle_rsc_0_0_i_bcwt_drv <= '0';
      ELSE
        twiddle_rsc_0_0_i_bcwt_drv <= NOT((NOT(twiddle_rsc_0_0_i_bcwt_drv OR twiddle_rsc_0_0_i_biwt))
            OR twiddle_rsc_0_0_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( twiddle_rsc_0_0_i_biwt = '1' ) THEN
        twiddle_rsc_0_0_i_s_din_bfwt <= twiddle_rsc_0_0_i_s_din;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_0_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_0_i_biwt : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_bdwt : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_bcwt : IN STD_LOGIC;
    twiddle_rsc_0_0_i_s_re_core_sct : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_s_rrdy : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_0_i_ogwt : STD_LOGIC;

BEGIN
  twiddle_rsc_0_0_i_bdwt <= twiddle_rsc_0_0_i_oswt AND core_wen;
  twiddle_rsc_0_0_i_biwt <= twiddle_rsc_0_0_i_ogwt AND twiddle_rsc_0_0_i_s_rrdy;
  twiddle_rsc_0_0_i_ogwt <= twiddle_rsc_0_0_i_oswt AND (NOT twiddle_rsc_0_0_i_bcwt);
  twiddle_rsc_0_0_i_s_re_core_sct <= twiddle_rsc_0_0_i_ogwt;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_31_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_31_i_biwt : IN STD_LOGIC;
    xt_rsc_1_31_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_31_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_31_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_31_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_31_i_qa_d, xt_rsc_1_31_i_qa_d_bfwt,
      xt_rsc_1_31_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_31_i_bcwt <= '0';
      ELSE
        xt_rsc_1_31_i_bcwt <= NOT((NOT(xt_rsc_1_31_i_bcwt OR xt_rsc_1_31_i_biwt))
            OR xt_rsc_1_31_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_31_i_biwt = '1' ) THEN
        xt_rsc_1_31_i_qa_d_bfwt <= xt_rsc_1_31_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_31_i_oswt : IN STD_LOGIC;
    xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_31_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_31_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_31_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_31_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_31_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_31_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_31_i_bdwt <= xt_rsc_1_31_i_oswt AND core_wen;
  xt_rsc_1_31_i_biwt <= (NOT core_wten) AND xt_rsc_1_31_i_oswt;
  xt_rsc_1_31_i_wea_d_core_sct_pff <= xt_rsc_1_31_i_wea_d_core_psct_pff AND xt_rsc_1_31_i_dswt_pff;
  xt_rsc_1_31_i_dswt_pff <= core_wen AND xt_rsc_1_31_i_oswt_pff;
  xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_31_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_30_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_30_i_biwt : IN STD_LOGIC;
    xt_rsc_1_30_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_30_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_30_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_30_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_30_i_qa_d, xt_rsc_1_30_i_qa_d_bfwt,
      xt_rsc_1_30_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_30_i_bcwt <= '0';
      ELSE
        xt_rsc_1_30_i_bcwt <= NOT((NOT(xt_rsc_1_30_i_bcwt OR xt_rsc_1_30_i_biwt))
            OR xt_rsc_1_30_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_30_i_biwt = '1' ) THEN
        xt_rsc_1_30_i_qa_d_bfwt <= xt_rsc_1_30_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_30_i_oswt : IN STD_LOGIC;
    xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_30_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_30_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_30_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_30_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_30_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_30_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_30_i_bdwt <= xt_rsc_1_30_i_oswt AND core_wen;
  xt_rsc_1_30_i_biwt <= (NOT core_wten) AND xt_rsc_1_30_i_oswt;
  xt_rsc_1_30_i_wea_d_core_sct_pff <= xt_rsc_1_30_i_wea_d_core_psct_pff AND xt_rsc_1_30_i_dswt_pff;
  xt_rsc_1_30_i_dswt_pff <= core_wen AND xt_rsc_1_30_i_oswt_pff;
  xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_30_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_29_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_29_i_biwt : IN STD_LOGIC;
    xt_rsc_1_29_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_29_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_29_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_29_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_29_i_qa_d, xt_rsc_1_29_i_qa_d_bfwt,
      xt_rsc_1_29_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_29_i_bcwt <= '0';
      ELSE
        xt_rsc_1_29_i_bcwt <= NOT((NOT(xt_rsc_1_29_i_bcwt OR xt_rsc_1_29_i_biwt))
            OR xt_rsc_1_29_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_29_i_biwt = '1' ) THEN
        xt_rsc_1_29_i_qa_d_bfwt <= xt_rsc_1_29_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_29_i_oswt : IN STD_LOGIC;
    xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_29_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_29_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_29_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_29_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_29_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_29_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_29_i_bdwt <= xt_rsc_1_29_i_oswt AND core_wen;
  xt_rsc_1_29_i_biwt <= (NOT core_wten) AND xt_rsc_1_29_i_oswt;
  xt_rsc_1_29_i_wea_d_core_sct_pff <= xt_rsc_1_29_i_wea_d_core_psct_pff AND xt_rsc_1_29_i_dswt_pff;
  xt_rsc_1_29_i_dswt_pff <= core_wen AND xt_rsc_1_29_i_oswt_pff;
  xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_29_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_28_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_28_i_biwt : IN STD_LOGIC;
    xt_rsc_1_28_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_28_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_28_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_28_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_28_i_qa_d, xt_rsc_1_28_i_qa_d_bfwt,
      xt_rsc_1_28_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_28_i_bcwt <= '0';
      ELSE
        xt_rsc_1_28_i_bcwt <= NOT((NOT(xt_rsc_1_28_i_bcwt OR xt_rsc_1_28_i_biwt))
            OR xt_rsc_1_28_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_28_i_biwt = '1' ) THEN
        xt_rsc_1_28_i_qa_d_bfwt <= xt_rsc_1_28_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_28_i_oswt : IN STD_LOGIC;
    xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_28_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_28_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_28_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_28_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_28_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_28_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_28_i_bdwt <= xt_rsc_1_28_i_oswt AND core_wen;
  xt_rsc_1_28_i_biwt <= (NOT core_wten) AND xt_rsc_1_28_i_oswt;
  xt_rsc_1_28_i_wea_d_core_sct_pff <= xt_rsc_1_28_i_wea_d_core_psct_pff AND xt_rsc_1_28_i_dswt_pff;
  xt_rsc_1_28_i_dswt_pff <= core_wen AND xt_rsc_1_28_i_oswt_pff;
  xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_28_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_27_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_27_i_biwt : IN STD_LOGIC;
    xt_rsc_1_27_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_27_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_27_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_27_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_27_i_qa_d, xt_rsc_1_27_i_qa_d_bfwt,
      xt_rsc_1_27_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_27_i_bcwt <= '0';
      ELSE
        xt_rsc_1_27_i_bcwt <= NOT((NOT(xt_rsc_1_27_i_bcwt OR xt_rsc_1_27_i_biwt))
            OR xt_rsc_1_27_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_27_i_biwt = '1' ) THEN
        xt_rsc_1_27_i_qa_d_bfwt <= xt_rsc_1_27_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_27_i_oswt : IN STD_LOGIC;
    xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_27_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_27_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_27_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_27_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_27_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_27_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_27_i_bdwt <= xt_rsc_1_27_i_oswt AND core_wen;
  xt_rsc_1_27_i_biwt <= (NOT core_wten) AND xt_rsc_1_27_i_oswt;
  xt_rsc_1_27_i_wea_d_core_sct_pff <= xt_rsc_1_27_i_wea_d_core_psct_pff AND xt_rsc_1_27_i_dswt_pff;
  xt_rsc_1_27_i_dswt_pff <= core_wen AND xt_rsc_1_27_i_oswt_pff;
  xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_27_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_26_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_26_i_biwt : IN STD_LOGIC;
    xt_rsc_1_26_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_26_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_26_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_26_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_26_i_qa_d, xt_rsc_1_26_i_qa_d_bfwt,
      xt_rsc_1_26_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_26_i_bcwt <= '0';
      ELSE
        xt_rsc_1_26_i_bcwt <= NOT((NOT(xt_rsc_1_26_i_bcwt OR xt_rsc_1_26_i_biwt))
            OR xt_rsc_1_26_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_26_i_biwt = '1' ) THEN
        xt_rsc_1_26_i_qa_d_bfwt <= xt_rsc_1_26_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_26_i_oswt : IN STD_LOGIC;
    xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_26_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_26_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_26_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_26_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_26_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_26_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_26_i_bdwt <= xt_rsc_1_26_i_oswt AND core_wen;
  xt_rsc_1_26_i_biwt <= (NOT core_wten) AND xt_rsc_1_26_i_oswt;
  xt_rsc_1_26_i_wea_d_core_sct_pff <= xt_rsc_1_26_i_wea_d_core_psct_pff AND xt_rsc_1_26_i_dswt_pff;
  xt_rsc_1_26_i_dswt_pff <= core_wen AND xt_rsc_1_26_i_oswt_pff;
  xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_26_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_25_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_25_i_biwt : IN STD_LOGIC;
    xt_rsc_1_25_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_25_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_25_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_25_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_25_i_qa_d, xt_rsc_1_25_i_qa_d_bfwt,
      xt_rsc_1_25_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_25_i_bcwt <= '0';
      ELSE
        xt_rsc_1_25_i_bcwt <= NOT((NOT(xt_rsc_1_25_i_bcwt OR xt_rsc_1_25_i_biwt))
            OR xt_rsc_1_25_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_25_i_biwt = '1' ) THEN
        xt_rsc_1_25_i_qa_d_bfwt <= xt_rsc_1_25_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_25_i_oswt : IN STD_LOGIC;
    xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_25_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_25_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_25_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_25_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_25_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_25_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_25_i_bdwt <= xt_rsc_1_25_i_oswt AND core_wen;
  xt_rsc_1_25_i_biwt <= (NOT core_wten) AND xt_rsc_1_25_i_oswt;
  xt_rsc_1_25_i_wea_d_core_sct_pff <= xt_rsc_1_25_i_wea_d_core_psct_pff AND xt_rsc_1_25_i_dswt_pff;
  xt_rsc_1_25_i_dswt_pff <= core_wen AND xt_rsc_1_25_i_oswt_pff;
  xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_25_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_24_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_24_i_biwt : IN STD_LOGIC;
    xt_rsc_1_24_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_24_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_24_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_24_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_24_i_qa_d, xt_rsc_1_24_i_qa_d_bfwt,
      xt_rsc_1_24_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_24_i_bcwt <= '0';
      ELSE
        xt_rsc_1_24_i_bcwt <= NOT((NOT(xt_rsc_1_24_i_bcwt OR xt_rsc_1_24_i_biwt))
            OR xt_rsc_1_24_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_24_i_biwt = '1' ) THEN
        xt_rsc_1_24_i_qa_d_bfwt <= xt_rsc_1_24_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_24_i_oswt : IN STD_LOGIC;
    xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_24_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_24_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_24_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_24_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_24_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_24_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_24_i_bdwt <= xt_rsc_1_24_i_oswt AND core_wen;
  xt_rsc_1_24_i_biwt <= (NOT core_wten) AND xt_rsc_1_24_i_oswt;
  xt_rsc_1_24_i_wea_d_core_sct_pff <= xt_rsc_1_24_i_wea_d_core_psct_pff AND xt_rsc_1_24_i_dswt_pff;
  xt_rsc_1_24_i_dswt_pff <= core_wen AND xt_rsc_1_24_i_oswt_pff;
  xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_24_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_23_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_23_i_biwt : IN STD_LOGIC;
    xt_rsc_1_23_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_23_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_23_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_23_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_23_i_qa_d, xt_rsc_1_23_i_qa_d_bfwt,
      xt_rsc_1_23_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_23_i_bcwt <= '0';
      ELSE
        xt_rsc_1_23_i_bcwt <= NOT((NOT(xt_rsc_1_23_i_bcwt OR xt_rsc_1_23_i_biwt))
            OR xt_rsc_1_23_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_23_i_biwt = '1' ) THEN
        xt_rsc_1_23_i_qa_d_bfwt <= xt_rsc_1_23_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_23_i_oswt : IN STD_LOGIC;
    xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_23_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_23_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_23_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_23_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_23_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_23_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_23_i_bdwt <= xt_rsc_1_23_i_oswt AND core_wen;
  xt_rsc_1_23_i_biwt <= (NOT core_wten) AND xt_rsc_1_23_i_oswt;
  xt_rsc_1_23_i_wea_d_core_sct_pff <= xt_rsc_1_23_i_wea_d_core_psct_pff AND xt_rsc_1_23_i_dswt_pff;
  xt_rsc_1_23_i_dswt_pff <= core_wen AND xt_rsc_1_23_i_oswt_pff;
  xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_23_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_22_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_22_i_biwt : IN STD_LOGIC;
    xt_rsc_1_22_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_22_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_22_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_22_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_22_i_qa_d, xt_rsc_1_22_i_qa_d_bfwt,
      xt_rsc_1_22_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_22_i_bcwt <= '0';
      ELSE
        xt_rsc_1_22_i_bcwt <= NOT((NOT(xt_rsc_1_22_i_bcwt OR xt_rsc_1_22_i_biwt))
            OR xt_rsc_1_22_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_22_i_biwt = '1' ) THEN
        xt_rsc_1_22_i_qa_d_bfwt <= xt_rsc_1_22_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_22_i_oswt : IN STD_LOGIC;
    xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_22_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_22_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_22_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_22_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_22_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_22_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_22_i_bdwt <= xt_rsc_1_22_i_oswt AND core_wen;
  xt_rsc_1_22_i_biwt <= (NOT core_wten) AND xt_rsc_1_22_i_oswt;
  xt_rsc_1_22_i_wea_d_core_sct_pff <= xt_rsc_1_22_i_wea_d_core_psct_pff AND xt_rsc_1_22_i_dswt_pff;
  xt_rsc_1_22_i_dswt_pff <= core_wen AND xt_rsc_1_22_i_oswt_pff;
  xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_22_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_21_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_21_i_biwt : IN STD_LOGIC;
    xt_rsc_1_21_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_21_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_21_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_21_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_21_i_qa_d, xt_rsc_1_21_i_qa_d_bfwt,
      xt_rsc_1_21_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_21_i_bcwt <= '0';
      ELSE
        xt_rsc_1_21_i_bcwt <= NOT((NOT(xt_rsc_1_21_i_bcwt OR xt_rsc_1_21_i_biwt))
            OR xt_rsc_1_21_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_21_i_biwt = '1' ) THEN
        xt_rsc_1_21_i_qa_d_bfwt <= xt_rsc_1_21_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_21_i_oswt : IN STD_LOGIC;
    xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_21_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_21_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_21_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_21_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_21_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_21_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_21_i_bdwt <= xt_rsc_1_21_i_oswt AND core_wen;
  xt_rsc_1_21_i_biwt <= (NOT core_wten) AND xt_rsc_1_21_i_oswt;
  xt_rsc_1_21_i_wea_d_core_sct_pff <= xt_rsc_1_21_i_wea_d_core_psct_pff AND xt_rsc_1_21_i_dswt_pff;
  xt_rsc_1_21_i_dswt_pff <= core_wen AND xt_rsc_1_21_i_oswt_pff;
  xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_21_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_20_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_20_i_biwt : IN STD_LOGIC;
    xt_rsc_1_20_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_20_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_20_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_20_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_20_i_qa_d, xt_rsc_1_20_i_qa_d_bfwt,
      xt_rsc_1_20_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_20_i_bcwt <= '0';
      ELSE
        xt_rsc_1_20_i_bcwt <= NOT((NOT(xt_rsc_1_20_i_bcwt OR xt_rsc_1_20_i_biwt))
            OR xt_rsc_1_20_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_20_i_biwt = '1' ) THEN
        xt_rsc_1_20_i_qa_d_bfwt <= xt_rsc_1_20_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_20_i_oswt : IN STD_LOGIC;
    xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_20_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_20_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_20_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_20_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_20_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_20_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_20_i_bdwt <= xt_rsc_1_20_i_oswt AND core_wen;
  xt_rsc_1_20_i_biwt <= (NOT core_wten) AND xt_rsc_1_20_i_oswt;
  xt_rsc_1_20_i_wea_d_core_sct_pff <= xt_rsc_1_20_i_wea_d_core_psct_pff AND xt_rsc_1_20_i_dswt_pff;
  xt_rsc_1_20_i_dswt_pff <= core_wen AND xt_rsc_1_20_i_oswt_pff;
  xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_20_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_19_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_19_i_biwt : IN STD_LOGIC;
    xt_rsc_1_19_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_19_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_19_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_19_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_19_i_qa_d, xt_rsc_1_19_i_qa_d_bfwt,
      xt_rsc_1_19_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_19_i_bcwt <= '0';
      ELSE
        xt_rsc_1_19_i_bcwt <= NOT((NOT(xt_rsc_1_19_i_bcwt OR xt_rsc_1_19_i_biwt))
            OR xt_rsc_1_19_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_19_i_biwt = '1' ) THEN
        xt_rsc_1_19_i_qa_d_bfwt <= xt_rsc_1_19_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_19_i_oswt : IN STD_LOGIC;
    xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_19_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_19_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_19_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_19_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_19_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_19_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_19_i_bdwt <= xt_rsc_1_19_i_oswt AND core_wen;
  xt_rsc_1_19_i_biwt <= (NOT core_wten) AND xt_rsc_1_19_i_oswt;
  xt_rsc_1_19_i_wea_d_core_sct_pff <= xt_rsc_1_19_i_wea_d_core_psct_pff AND xt_rsc_1_19_i_dswt_pff;
  xt_rsc_1_19_i_dswt_pff <= core_wen AND xt_rsc_1_19_i_oswt_pff;
  xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_19_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_18_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_18_i_biwt : IN STD_LOGIC;
    xt_rsc_1_18_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_18_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_18_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_18_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_18_i_qa_d, xt_rsc_1_18_i_qa_d_bfwt,
      xt_rsc_1_18_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_18_i_bcwt <= '0';
      ELSE
        xt_rsc_1_18_i_bcwt <= NOT((NOT(xt_rsc_1_18_i_bcwt OR xt_rsc_1_18_i_biwt))
            OR xt_rsc_1_18_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_18_i_biwt = '1' ) THEN
        xt_rsc_1_18_i_qa_d_bfwt <= xt_rsc_1_18_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_18_i_oswt : IN STD_LOGIC;
    xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_18_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_18_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_18_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_18_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_18_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_18_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_18_i_bdwt <= xt_rsc_1_18_i_oswt AND core_wen;
  xt_rsc_1_18_i_biwt <= (NOT core_wten) AND xt_rsc_1_18_i_oswt;
  xt_rsc_1_18_i_wea_d_core_sct_pff <= xt_rsc_1_18_i_wea_d_core_psct_pff AND xt_rsc_1_18_i_dswt_pff;
  xt_rsc_1_18_i_dswt_pff <= core_wen AND xt_rsc_1_18_i_oswt_pff;
  xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_18_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_17_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_17_i_biwt : IN STD_LOGIC;
    xt_rsc_1_17_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_17_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_17_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_17_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_17_i_qa_d, xt_rsc_1_17_i_qa_d_bfwt,
      xt_rsc_1_17_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_17_i_bcwt <= '0';
      ELSE
        xt_rsc_1_17_i_bcwt <= NOT((NOT(xt_rsc_1_17_i_bcwt OR xt_rsc_1_17_i_biwt))
            OR xt_rsc_1_17_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_17_i_biwt = '1' ) THEN
        xt_rsc_1_17_i_qa_d_bfwt <= xt_rsc_1_17_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_17_i_oswt : IN STD_LOGIC;
    xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_17_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_17_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_17_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_17_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_17_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_17_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_17_i_bdwt <= xt_rsc_1_17_i_oswt AND core_wen;
  xt_rsc_1_17_i_biwt <= (NOT core_wten) AND xt_rsc_1_17_i_oswt;
  xt_rsc_1_17_i_wea_d_core_sct_pff <= xt_rsc_1_17_i_wea_d_core_psct_pff AND xt_rsc_1_17_i_dswt_pff;
  xt_rsc_1_17_i_dswt_pff <= core_wen AND xt_rsc_1_17_i_oswt_pff;
  xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_17_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_16_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_16_i_biwt : IN STD_LOGIC;
    xt_rsc_1_16_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_16_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_16_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_16_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_16_i_qa_d, xt_rsc_1_16_i_qa_d_bfwt,
      xt_rsc_1_16_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_16_i_bcwt <= '0';
      ELSE
        xt_rsc_1_16_i_bcwt <= NOT((NOT(xt_rsc_1_16_i_bcwt OR xt_rsc_1_16_i_biwt))
            OR xt_rsc_1_16_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_16_i_biwt = '1' ) THEN
        xt_rsc_1_16_i_qa_d_bfwt <= xt_rsc_1_16_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_16_i_oswt : IN STD_LOGIC;
    xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_16_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_16_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_16_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_16_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_16_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_16_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_16_i_bdwt <= xt_rsc_1_16_i_oswt AND core_wen;
  xt_rsc_1_16_i_biwt <= (NOT core_wten) AND xt_rsc_1_16_i_oswt;
  xt_rsc_1_16_i_wea_d_core_sct_pff <= xt_rsc_1_16_i_wea_d_core_psct_pff AND xt_rsc_1_16_i_dswt_pff;
  xt_rsc_1_16_i_dswt_pff <= core_wen AND xt_rsc_1_16_i_oswt_pff;
  xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_16_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_15_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_15_i_biwt : IN STD_LOGIC;
    xt_rsc_1_15_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_15_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_15_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_15_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_15_i_qa_d, xt_rsc_1_15_i_qa_d_bfwt,
      xt_rsc_1_15_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_15_i_bcwt <= '0';
      ELSE
        xt_rsc_1_15_i_bcwt <= NOT((NOT(xt_rsc_1_15_i_bcwt OR xt_rsc_1_15_i_biwt))
            OR xt_rsc_1_15_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_15_i_biwt = '1' ) THEN
        xt_rsc_1_15_i_qa_d_bfwt <= xt_rsc_1_15_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_15_i_oswt : IN STD_LOGIC;
    xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_15_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_15_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_15_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_15_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_15_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_15_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_15_i_bdwt <= xt_rsc_1_15_i_oswt AND core_wen;
  xt_rsc_1_15_i_biwt <= (NOT core_wten) AND xt_rsc_1_15_i_oswt;
  xt_rsc_1_15_i_wea_d_core_sct_pff <= xt_rsc_1_15_i_wea_d_core_psct_pff AND xt_rsc_1_15_i_dswt_pff;
  xt_rsc_1_15_i_dswt_pff <= core_wen AND xt_rsc_1_15_i_oswt_pff;
  xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_15_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_14_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_14_i_biwt : IN STD_LOGIC;
    xt_rsc_1_14_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_14_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_14_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_14_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_14_i_qa_d, xt_rsc_1_14_i_qa_d_bfwt,
      xt_rsc_1_14_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_14_i_bcwt <= '0';
      ELSE
        xt_rsc_1_14_i_bcwt <= NOT((NOT(xt_rsc_1_14_i_bcwt OR xt_rsc_1_14_i_biwt))
            OR xt_rsc_1_14_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_14_i_biwt = '1' ) THEN
        xt_rsc_1_14_i_qa_d_bfwt <= xt_rsc_1_14_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_14_i_oswt : IN STD_LOGIC;
    xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_14_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_14_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_14_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_14_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_14_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_14_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_14_i_bdwt <= xt_rsc_1_14_i_oswt AND core_wen;
  xt_rsc_1_14_i_biwt <= (NOT core_wten) AND xt_rsc_1_14_i_oswt;
  xt_rsc_1_14_i_wea_d_core_sct_pff <= xt_rsc_1_14_i_wea_d_core_psct_pff AND xt_rsc_1_14_i_dswt_pff;
  xt_rsc_1_14_i_dswt_pff <= core_wen AND xt_rsc_1_14_i_oswt_pff;
  xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_14_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_13_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_13_i_biwt : IN STD_LOGIC;
    xt_rsc_1_13_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_13_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_13_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_13_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_13_i_qa_d, xt_rsc_1_13_i_qa_d_bfwt,
      xt_rsc_1_13_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_13_i_bcwt <= '0';
      ELSE
        xt_rsc_1_13_i_bcwt <= NOT((NOT(xt_rsc_1_13_i_bcwt OR xt_rsc_1_13_i_biwt))
            OR xt_rsc_1_13_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_13_i_biwt = '1' ) THEN
        xt_rsc_1_13_i_qa_d_bfwt <= xt_rsc_1_13_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_13_i_oswt : IN STD_LOGIC;
    xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_13_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_13_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_13_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_13_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_13_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_13_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_13_i_bdwt <= xt_rsc_1_13_i_oswt AND core_wen;
  xt_rsc_1_13_i_biwt <= (NOT core_wten) AND xt_rsc_1_13_i_oswt;
  xt_rsc_1_13_i_wea_d_core_sct_pff <= xt_rsc_1_13_i_wea_d_core_psct_pff AND xt_rsc_1_13_i_dswt_pff;
  xt_rsc_1_13_i_dswt_pff <= core_wen AND xt_rsc_1_13_i_oswt_pff;
  xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_13_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_12_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_12_i_biwt : IN STD_LOGIC;
    xt_rsc_1_12_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_12_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_12_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_12_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_12_i_qa_d, xt_rsc_1_12_i_qa_d_bfwt,
      xt_rsc_1_12_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_12_i_bcwt <= '0';
      ELSE
        xt_rsc_1_12_i_bcwt <= NOT((NOT(xt_rsc_1_12_i_bcwt OR xt_rsc_1_12_i_biwt))
            OR xt_rsc_1_12_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_12_i_biwt = '1' ) THEN
        xt_rsc_1_12_i_qa_d_bfwt <= xt_rsc_1_12_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_12_i_oswt : IN STD_LOGIC;
    xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_12_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_12_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_12_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_12_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_12_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_12_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_12_i_bdwt <= xt_rsc_1_12_i_oswt AND core_wen;
  xt_rsc_1_12_i_biwt <= (NOT core_wten) AND xt_rsc_1_12_i_oswt;
  xt_rsc_1_12_i_wea_d_core_sct_pff <= xt_rsc_1_12_i_wea_d_core_psct_pff AND xt_rsc_1_12_i_dswt_pff;
  xt_rsc_1_12_i_dswt_pff <= core_wen AND xt_rsc_1_12_i_oswt_pff;
  xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_12_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_11_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_11_i_biwt : IN STD_LOGIC;
    xt_rsc_1_11_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_11_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_11_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_11_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_11_i_qa_d, xt_rsc_1_11_i_qa_d_bfwt,
      xt_rsc_1_11_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_11_i_bcwt <= '0';
      ELSE
        xt_rsc_1_11_i_bcwt <= NOT((NOT(xt_rsc_1_11_i_bcwt OR xt_rsc_1_11_i_biwt))
            OR xt_rsc_1_11_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_11_i_biwt = '1' ) THEN
        xt_rsc_1_11_i_qa_d_bfwt <= xt_rsc_1_11_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_11_i_oswt : IN STD_LOGIC;
    xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_11_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_11_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_11_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_11_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_11_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_11_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_11_i_bdwt <= xt_rsc_1_11_i_oswt AND core_wen;
  xt_rsc_1_11_i_biwt <= (NOT core_wten) AND xt_rsc_1_11_i_oswt;
  xt_rsc_1_11_i_wea_d_core_sct_pff <= xt_rsc_1_11_i_wea_d_core_psct_pff AND xt_rsc_1_11_i_dswt_pff;
  xt_rsc_1_11_i_dswt_pff <= core_wen AND xt_rsc_1_11_i_oswt_pff;
  xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_11_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_10_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_10_i_biwt : IN STD_LOGIC;
    xt_rsc_1_10_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_10_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_10_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_10_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_10_i_qa_d, xt_rsc_1_10_i_qa_d_bfwt,
      xt_rsc_1_10_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_10_i_bcwt <= '0';
      ELSE
        xt_rsc_1_10_i_bcwt <= NOT((NOT(xt_rsc_1_10_i_bcwt OR xt_rsc_1_10_i_biwt))
            OR xt_rsc_1_10_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_10_i_biwt = '1' ) THEN
        xt_rsc_1_10_i_qa_d_bfwt <= xt_rsc_1_10_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_10_i_oswt : IN STD_LOGIC;
    xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_10_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_10_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_10_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_10_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_10_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_10_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_10_i_bdwt <= xt_rsc_1_10_i_oswt AND core_wen;
  xt_rsc_1_10_i_biwt <= (NOT core_wten) AND xt_rsc_1_10_i_oswt;
  xt_rsc_1_10_i_wea_d_core_sct_pff <= xt_rsc_1_10_i_wea_d_core_psct_pff AND xt_rsc_1_10_i_dswt_pff;
  xt_rsc_1_10_i_dswt_pff <= core_wen AND xt_rsc_1_10_i_oswt_pff;
  xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_10_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_9_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_9_i_biwt : IN STD_LOGIC;
    xt_rsc_1_9_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_9_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_9_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_9_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_9_i_qa_d, xt_rsc_1_9_i_qa_d_bfwt,
      xt_rsc_1_9_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_9_i_bcwt <= '0';
      ELSE
        xt_rsc_1_9_i_bcwt <= NOT((NOT(xt_rsc_1_9_i_bcwt OR xt_rsc_1_9_i_biwt)) OR
            xt_rsc_1_9_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_9_i_biwt = '1' ) THEN
        xt_rsc_1_9_i_qa_d_bfwt <= xt_rsc_1_9_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_9_i_oswt : IN STD_LOGIC;
    xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_9_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_9_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_9_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_9_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_9_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_9_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_9_i_bdwt <= xt_rsc_1_9_i_oswt AND core_wen;
  xt_rsc_1_9_i_biwt <= (NOT core_wten) AND xt_rsc_1_9_i_oswt;
  xt_rsc_1_9_i_wea_d_core_sct_pff <= xt_rsc_1_9_i_wea_d_core_psct_pff AND xt_rsc_1_9_i_dswt_pff;
  xt_rsc_1_9_i_dswt_pff <= core_wen AND xt_rsc_1_9_i_oswt_pff;
  xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_9_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_8_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_8_i_biwt : IN STD_LOGIC;
    xt_rsc_1_8_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_8_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_8_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_8_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_8_i_qa_d, xt_rsc_1_8_i_qa_d_bfwt,
      xt_rsc_1_8_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_8_i_bcwt <= '0';
      ELSE
        xt_rsc_1_8_i_bcwt <= NOT((NOT(xt_rsc_1_8_i_bcwt OR xt_rsc_1_8_i_biwt)) OR
            xt_rsc_1_8_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_8_i_biwt = '1' ) THEN
        xt_rsc_1_8_i_qa_d_bfwt <= xt_rsc_1_8_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_8_i_oswt : IN STD_LOGIC;
    xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_8_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_8_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_8_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_8_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_8_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_8_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_8_i_bdwt <= xt_rsc_1_8_i_oswt AND core_wen;
  xt_rsc_1_8_i_biwt <= (NOT core_wten) AND xt_rsc_1_8_i_oswt;
  xt_rsc_1_8_i_wea_d_core_sct_pff <= xt_rsc_1_8_i_wea_d_core_psct_pff AND xt_rsc_1_8_i_dswt_pff;
  xt_rsc_1_8_i_dswt_pff <= core_wen AND xt_rsc_1_8_i_oswt_pff;
  xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_8_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_7_i_biwt : IN STD_LOGIC;
    xt_rsc_1_7_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_7_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_7_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_7_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_7_i_qa_d, xt_rsc_1_7_i_qa_d_bfwt,
      xt_rsc_1_7_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_7_i_bcwt <= '0';
      ELSE
        xt_rsc_1_7_i_bcwt <= NOT((NOT(xt_rsc_1_7_i_bcwt OR xt_rsc_1_7_i_biwt)) OR
            xt_rsc_1_7_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_7_i_biwt = '1' ) THEN
        xt_rsc_1_7_i_qa_d_bfwt <= xt_rsc_1_7_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_7_i_oswt : IN STD_LOGIC;
    xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_7_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_7_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_7_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_7_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_7_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_7_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_7_i_bdwt <= xt_rsc_1_7_i_oswt AND core_wen;
  xt_rsc_1_7_i_biwt <= (NOT core_wten) AND xt_rsc_1_7_i_oswt;
  xt_rsc_1_7_i_wea_d_core_sct_pff <= xt_rsc_1_7_i_wea_d_core_psct_pff AND xt_rsc_1_7_i_dswt_pff;
  xt_rsc_1_7_i_dswt_pff <= core_wen AND xt_rsc_1_7_i_oswt_pff;
  xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_7_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_6_i_biwt : IN STD_LOGIC;
    xt_rsc_1_6_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_6_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_6_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_6_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_6_i_qa_d, xt_rsc_1_6_i_qa_d_bfwt,
      xt_rsc_1_6_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_6_i_bcwt <= '0';
      ELSE
        xt_rsc_1_6_i_bcwt <= NOT((NOT(xt_rsc_1_6_i_bcwt OR xt_rsc_1_6_i_biwt)) OR
            xt_rsc_1_6_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_6_i_biwt = '1' ) THEN
        xt_rsc_1_6_i_qa_d_bfwt <= xt_rsc_1_6_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_6_i_oswt : IN STD_LOGIC;
    xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_6_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_6_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_6_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_6_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_6_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_6_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_6_i_bdwt <= xt_rsc_1_6_i_oswt AND core_wen;
  xt_rsc_1_6_i_biwt <= (NOT core_wten) AND xt_rsc_1_6_i_oswt;
  xt_rsc_1_6_i_wea_d_core_sct_pff <= xt_rsc_1_6_i_wea_d_core_psct_pff AND xt_rsc_1_6_i_dswt_pff;
  xt_rsc_1_6_i_dswt_pff <= core_wen AND xt_rsc_1_6_i_oswt_pff;
  xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_6_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_5_i_biwt : IN STD_LOGIC;
    xt_rsc_1_5_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_5_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_5_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_5_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_5_i_qa_d, xt_rsc_1_5_i_qa_d_bfwt,
      xt_rsc_1_5_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_5_i_bcwt <= '0';
      ELSE
        xt_rsc_1_5_i_bcwt <= NOT((NOT(xt_rsc_1_5_i_bcwt OR xt_rsc_1_5_i_biwt)) OR
            xt_rsc_1_5_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_5_i_biwt = '1' ) THEN
        xt_rsc_1_5_i_qa_d_bfwt <= xt_rsc_1_5_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_5_i_oswt : IN STD_LOGIC;
    xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_5_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_5_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_5_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_5_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_5_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_5_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_5_i_bdwt <= xt_rsc_1_5_i_oswt AND core_wen;
  xt_rsc_1_5_i_biwt <= (NOT core_wten) AND xt_rsc_1_5_i_oswt;
  xt_rsc_1_5_i_wea_d_core_sct_pff <= xt_rsc_1_5_i_wea_d_core_psct_pff AND xt_rsc_1_5_i_dswt_pff;
  xt_rsc_1_5_i_dswt_pff <= core_wen AND xt_rsc_1_5_i_oswt_pff;
  xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_5_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_4_i_biwt : IN STD_LOGIC;
    xt_rsc_1_4_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_4_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_4_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_4_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_4_i_qa_d, xt_rsc_1_4_i_qa_d_bfwt,
      xt_rsc_1_4_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_4_i_bcwt <= '0';
      ELSE
        xt_rsc_1_4_i_bcwt <= NOT((NOT(xt_rsc_1_4_i_bcwt OR xt_rsc_1_4_i_biwt)) OR
            xt_rsc_1_4_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_4_i_biwt = '1' ) THEN
        xt_rsc_1_4_i_qa_d_bfwt <= xt_rsc_1_4_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_4_i_oswt : IN STD_LOGIC;
    xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_4_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_4_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_4_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_4_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_4_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_4_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_4_i_bdwt <= xt_rsc_1_4_i_oswt AND core_wen;
  xt_rsc_1_4_i_biwt <= (NOT core_wten) AND xt_rsc_1_4_i_oswt;
  xt_rsc_1_4_i_wea_d_core_sct_pff <= xt_rsc_1_4_i_wea_d_core_psct_pff AND xt_rsc_1_4_i_dswt_pff;
  xt_rsc_1_4_i_dswt_pff <= core_wen AND xt_rsc_1_4_i_oswt_pff;
  xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_4_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_3_i_biwt : IN STD_LOGIC;
    xt_rsc_1_3_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_3_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_3_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_3_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_3_i_qa_d, xt_rsc_1_3_i_qa_d_bfwt,
      xt_rsc_1_3_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_3_i_bcwt <= '0';
      ELSE
        xt_rsc_1_3_i_bcwt <= NOT((NOT(xt_rsc_1_3_i_bcwt OR xt_rsc_1_3_i_biwt)) OR
            xt_rsc_1_3_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_3_i_biwt = '1' ) THEN
        xt_rsc_1_3_i_qa_d_bfwt <= xt_rsc_1_3_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_3_i_oswt : IN STD_LOGIC;
    xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_3_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_3_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_3_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_3_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_3_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_3_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_3_i_bdwt <= xt_rsc_1_3_i_oswt AND core_wen;
  xt_rsc_1_3_i_biwt <= (NOT core_wten) AND xt_rsc_1_3_i_oswt;
  xt_rsc_1_3_i_wea_d_core_sct_pff <= xt_rsc_1_3_i_wea_d_core_psct_pff AND xt_rsc_1_3_i_dswt_pff;
  xt_rsc_1_3_i_dswt_pff <= core_wen AND xt_rsc_1_3_i_oswt_pff;
  xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_3_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_2_i_biwt : IN STD_LOGIC;
    xt_rsc_1_2_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_2_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_2_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_2_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_2_i_qa_d, xt_rsc_1_2_i_qa_d_bfwt,
      xt_rsc_1_2_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_2_i_bcwt <= '0';
      ELSE
        xt_rsc_1_2_i_bcwt <= NOT((NOT(xt_rsc_1_2_i_bcwt OR xt_rsc_1_2_i_biwt)) OR
            xt_rsc_1_2_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_2_i_biwt = '1' ) THEN
        xt_rsc_1_2_i_qa_d_bfwt <= xt_rsc_1_2_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_2_i_oswt : IN STD_LOGIC;
    xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_2_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_2_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_2_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_2_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_2_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_2_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_2_i_bdwt <= xt_rsc_1_2_i_oswt AND core_wen;
  xt_rsc_1_2_i_biwt <= (NOT core_wten) AND xt_rsc_1_2_i_oswt;
  xt_rsc_1_2_i_wea_d_core_sct_pff <= xt_rsc_1_2_i_wea_d_core_psct_pff AND xt_rsc_1_2_i_dswt_pff;
  xt_rsc_1_2_i_dswt_pff <= core_wen AND xt_rsc_1_2_i_oswt_pff;
  xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_2_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_1_i_biwt : IN STD_LOGIC;
    xt_rsc_1_1_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_1_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_1_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_1_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_1_i_qa_d, xt_rsc_1_1_i_qa_d_bfwt,
      xt_rsc_1_1_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_1_i_bcwt <= '0';
      ELSE
        xt_rsc_1_1_i_bcwt <= NOT((NOT(xt_rsc_1_1_i_bcwt OR xt_rsc_1_1_i_biwt)) OR
            xt_rsc_1_1_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_1_i_biwt = '1' ) THEN
        xt_rsc_1_1_i_qa_d_bfwt <= xt_rsc_1_1_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_1_i_oswt : IN STD_LOGIC;
    xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_1_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_1_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_1_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_1_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_1_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_1_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_1_i_bdwt <= xt_rsc_1_1_i_oswt AND core_wen;
  xt_rsc_1_1_i_biwt <= (NOT core_wten) AND xt_rsc_1_1_i_oswt;
  xt_rsc_1_1_i_wea_d_core_sct_pff <= xt_rsc_1_1_i_wea_d_core_psct_pff AND xt_rsc_1_1_i_dswt_pff;
  xt_rsc_1_1_i_dswt_pff <= core_wen AND xt_rsc_1_1_i_oswt_pff;
  xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_1_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_0_i_biwt : IN STD_LOGIC;
    xt_rsc_1_0_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_0_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_1_0_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_1_0_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_1_0_i_qa_d, xt_rsc_1_0_i_qa_d_bfwt,
      xt_rsc_1_0_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_1_0_i_bcwt <= '0';
      ELSE
        xt_rsc_1_0_i_bcwt <= NOT((NOT(xt_rsc_1_0_i_bcwt OR xt_rsc_1_0_i_biwt)) OR
            xt_rsc_1_0_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_1_0_i_biwt = '1' ) THEN
        xt_rsc_1_0_i_qa_d_bfwt <= xt_rsc_1_0_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_0_i_oswt : IN STD_LOGIC;
    xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_0_i_biwt : OUT STD_LOGIC;
    xt_rsc_1_0_i_bdwt : OUT STD_LOGIC;
    xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_1_0_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_1_0_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_0_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_0_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_1_0_i_bdwt <= xt_rsc_1_0_i_oswt AND core_wen;
  xt_rsc_1_0_i_biwt <= (NOT core_wten) AND xt_rsc_1_0_i_oswt;
  xt_rsc_1_0_i_wea_d_core_sct_pff <= xt_rsc_1_0_i_wea_d_core_psct_pff AND xt_rsc_1_0_i_dswt_pff;
  xt_rsc_1_0_i_dswt_pff <= core_wen AND xt_rsc_1_0_i_oswt_pff;
  xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_1_0_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_31_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_31_i_biwt : IN STD_LOGIC;
    xt_rsc_0_31_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_31_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_31_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_31_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_31_i_qa_d, xt_rsc_0_31_i_qa_d_bfwt,
      xt_rsc_0_31_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_31_i_bcwt <= '0';
      ELSE
        xt_rsc_0_31_i_bcwt <= NOT((NOT(xt_rsc_0_31_i_bcwt OR xt_rsc_0_31_i_biwt))
            OR xt_rsc_0_31_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_31_i_biwt = '1' ) THEN
        xt_rsc_0_31_i_qa_d_bfwt <= xt_rsc_0_31_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_31_i_oswt : IN STD_LOGIC;
    xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_31_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_31_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_31_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_31_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_31_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_31_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_31_i_bdwt <= xt_rsc_0_31_i_oswt AND core_wen;
  xt_rsc_0_31_i_biwt <= (NOT core_wten) AND xt_rsc_0_31_i_oswt;
  xt_rsc_0_31_i_wea_d_core_sct_pff <= xt_rsc_0_31_i_wea_d_core_psct_pff AND xt_rsc_0_31_i_dswt_pff;
  xt_rsc_0_31_i_dswt_pff <= core_wen AND xt_rsc_0_31_i_oswt_pff;
  xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_31_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_30_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_30_i_biwt : IN STD_LOGIC;
    xt_rsc_0_30_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_30_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_30_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_30_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_30_i_qa_d, xt_rsc_0_30_i_qa_d_bfwt,
      xt_rsc_0_30_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_30_i_bcwt <= '0';
      ELSE
        xt_rsc_0_30_i_bcwt <= NOT((NOT(xt_rsc_0_30_i_bcwt OR xt_rsc_0_30_i_biwt))
            OR xt_rsc_0_30_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_30_i_biwt = '1' ) THEN
        xt_rsc_0_30_i_qa_d_bfwt <= xt_rsc_0_30_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_30_i_oswt : IN STD_LOGIC;
    xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_30_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_30_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_30_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_30_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_30_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_30_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_30_i_bdwt <= xt_rsc_0_30_i_oswt AND core_wen;
  xt_rsc_0_30_i_biwt <= (NOT core_wten) AND xt_rsc_0_30_i_oswt;
  xt_rsc_0_30_i_wea_d_core_sct_pff <= xt_rsc_0_30_i_wea_d_core_psct_pff AND xt_rsc_0_30_i_dswt_pff;
  xt_rsc_0_30_i_dswt_pff <= core_wen AND xt_rsc_0_30_i_oswt_pff;
  xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_30_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_29_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_29_i_biwt : IN STD_LOGIC;
    xt_rsc_0_29_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_29_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_29_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_29_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_29_i_qa_d, xt_rsc_0_29_i_qa_d_bfwt,
      xt_rsc_0_29_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_29_i_bcwt <= '0';
      ELSE
        xt_rsc_0_29_i_bcwt <= NOT((NOT(xt_rsc_0_29_i_bcwt OR xt_rsc_0_29_i_biwt))
            OR xt_rsc_0_29_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_29_i_biwt = '1' ) THEN
        xt_rsc_0_29_i_qa_d_bfwt <= xt_rsc_0_29_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_29_i_oswt : IN STD_LOGIC;
    xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_29_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_29_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_29_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_29_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_29_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_29_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_29_i_bdwt <= xt_rsc_0_29_i_oswt AND core_wen;
  xt_rsc_0_29_i_biwt <= (NOT core_wten) AND xt_rsc_0_29_i_oswt;
  xt_rsc_0_29_i_wea_d_core_sct_pff <= xt_rsc_0_29_i_wea_d_core_psct_pff AND xt_rsc_0_29_i_dswt_pff;
  xt_rsc_0_29_i_dswt_pff <= core_wen AND xt_rsc_0_29_i_oswt_pff;
  xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_29_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_28_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_28_i_biwt : IN STD_LOGIC;
    xt_rsc_0_28_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_28_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_28_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_28_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_28_i_qa_d, xt_rsc_0_28_i_qa_d_bfwt,
      xt_rsc_0_28_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_28_i_bcwt <= '0';
      ELSE
        xt_rsc_0_28_i_bcwt <= NOT((NOT(xt_rsc_0_28_i_bcwt OR xt_rsc_0_28_i_biwt))
            OR xt_rsc_0_28_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_28_i_biwt = '1' ) THEN
        xt_rsc_0_28_i_qa_d_bfwt <= xt_rsc_0_28_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_28_i_oswt : IN STD_LOGIC;
    xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_28_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_28_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_28_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_28_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_28_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_28_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_28_i_bdwt <= xt_rsc_0_28_i_oswt AND core_wen;
  xt_rsc_0_28_i_biwt <= (NOT core_wten) AND xt_rsc_0_28_i_oswt;
  xt_rsc_0_28_i_wea_d_core_sct_pff <= xt_rsc_0_28_i_wea_d_core_psct_pff AND xt_rsc_0_28_i_dswt_pff;
  xt_rsc_0_28_i_dswt_pff <= core_wen AND xt_rsc_0_28_i_oswt_pff;
  xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_28_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_27_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_27_i_biwt : IN STD_LOGIC;
    xt_rsc_0_27_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_27_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_27_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_27_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_27_i_qa_d, xt_rsc_0_27_i_qa_d_bfwt,
      xt_rsc_0_27_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_27_i_bcwt <= '0';
      ELSE
        xt_rsc_0_27_i_bcwt <= NOT((NOT(xt_rsc_0_27_i_bcwt OR xt_rsc_0_27_i_biwt))
            OR xt_rsc_0_27_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_27_i_biwt = '1' ) THEN
        xt_rsc_0_27_i_qa_d_bfwt <= xt_rsc_0_27_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_27_i_oswt : IN STD_LOGIC;
    xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_27_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_27_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_27_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_27_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_27_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_27_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_27_i_bdwt <= xt_rsc_0_27_i_oswt AND core_wen;
  xt_rsc_0_27_i_biwt <= (NOT core_wten) AND xt_rsc_0_27_i_oswt;
  xt_rsc_0_27_i_wea_d_core_sct_pff <= xt_rsc_0_27_i_wea_d_core_psct_pff AND xt_rsc_0_27_i_dswt_pff;
  xt_rsc_0_27_i_dswt_pff <= core_wen AND xt_rsc_0_27_i_oswt_pff;
  xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_27_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_26_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_26_i_biwt : IN STD_LOGIC;
    xt_rsc_0_26_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_26_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_26_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_26_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_26_i_qa_d, xt_rsc_0_26_i_qa_d_bfwt,
      xt_rsc_0_26_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_26_i_bcwt <= '0';
      ELSE
        xt_rsc_0_26_i_bcwt <= NOT((NOT(xt_rsc_0_26_i_bcwt OR xt_rsc_0_26_i_biwt))
            OR xt_rsc_0_26_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_26_i_biwt = '1' ) THEN
        xt_rsc_0_26_i_qa_d_bfwt <= xt_rsc_0_26_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_26_i_oswt : IN STD_LOGIC;
    xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_26_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_26_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_26_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_26_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_26_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_26_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_26_i_bdwt <= xt_rsc_0_26_i_oswt AND core_wen;
  xt_rsc_0_26_i_biwt <= (NOT core_wten) AND xt_rsc_0_26_i_oswt;
  xt_rsc_0_26_i_wea_d_core_sct_pff <= xt_rsc_0_26_i_wea_d_core_psct_pff AND xt_rsc_0_26_i_dswt_pff;
  xt_rsc_0_26_i_dswt_pff <= core_wen AND xt_rsc_0_26_i_oswt_pff;
  xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_26_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_25_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_25_i_biwt : IN STD_LOGIC;
    xt_rsc_0_25_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_25_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_25_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_25_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_25_i_qa_d, xt_rsc_0_25_i_qa_d_bfwt,
      xt_rsc_0_25_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_25_i_bcwt <= '0';
      ELSE
        xt_rsc_0_25_i_bcwt <= NOT((NOT(xt_rsc_0_25_i_bcwt OR xt_rsc_0_25_i_biwt))
            OR xt_rsc_0_25_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_25_i_biwt = '1' ) THEN
        xt_rsc_0_25_i_qa_d_bfwt <= xt_rsc_0_25_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_25_i_oswt : IN STD_LOGIC;
    xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_25_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_25_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_25_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_25_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_25_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_25_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_25_i_bdwt <= xt_rsc_0_25_i_oswt AND core_wen;
  xt_rsc_0_25_i_biwt <= (NOT core_wten) AND xt_rsc_0_25_i_oswt;
  xt_rsc_0_25_i_wea_d_core_sct_pff <= xt_rsc_0_25_i_wea_d_core_psct_pff AND xt_rsc_0_25_i_dswt_pff;
  xt_rsc_0_25_i_dswt_pff <= core_wen AND xt_rsc_0_25_i_oswt_pff;
  xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_25_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_24_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_24_i_biwt : IN STD_LOGIC;
    xt_rsc_0_24_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_24_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_24_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_24_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_24_i_qa_d, xt_rsc_0_24_i_qa_d_bfwt,
      xt_rsc_0_24_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_24_i_bcwt <= '0';
      ELSE
        xt_rsc_0_24_i_bcwt <= NOT((NOT(xt_rsc_0_24_i_bcwt OR xt_rsc_0_24_i_biwt))
            OR xt_rsc_0_24_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_24_i_biwt = '1' ) THEN
        xt_rsc_0_24_i_qa_d_bfwt <= xt_rsc_0_24_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_24_i_oswt : IN STD_LOGIC;
    xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_24_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_24_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_24_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_24_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_24_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_24_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_24_i_bdwt <= xt_rsc_0_24_i_oswt AND core_wen;
  xt_rsc_0_24_i_biwt <= (NOT core_wten) AND xt_rsc_0_24_i_oswt;
  xt_rsc_0_24_i_wea_d_core_sct_pff <= xt_rsc_0_24_i_wea_d_core_psct_pff AND xt_rsc_0_24_i_dswt_pff;
  xt_rsc_0_24_i_dswt_pff <= core_wen AND xt_rsc_0_24_i_oswt_pff;
  xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_24_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_23_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_23_i_biwt : IN STD_LOGIC;
    xt_rsc_0_23_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_23_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_23_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_23_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_23_i_qa_d, xt_rsc_0_23_i_qa_d_bfwt,
      xt_rsc_0_23_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_23_i_bcwt <= '0';
      ELSE
        xt_rsc_0_23_i_bcwt <= NOT((NOT(xt_rsc_0_23_i_bcwt OR xt_rsc_0_23_i_biwt))
            OR xt_rsc_0_23_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_23_i_biwt = '1' ) THEN
        xt_rsc_0_23_i_qa_d_bfwt <= xt_rsc_0_23_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_23_i_oswt : IN STD_LOGIC;
    xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_23_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_23_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_23_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_23_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_23_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_23_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_23_i_bdwt <= xt_rsc_0_23_i_oswt AND core_wen;
  xt_rsc_0_23_i_biwt <= (NOT core_wten) AND xt_rsc_0_23_i_oswt;
  xt_rsc_0_23_i_wea_d_core_sct_pff <= xt_rsc_0_23_i_wea_d_core_psct_pff AND xt_rsc_0_23_i_dswt_pff;
  xt_rsc_0_23_i_dswt_pff <= core_wen AND xt_rsc_0_23_i_oswt_pff;
  xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_23_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_22_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_22_i_biwt : IN STD_LOGIC;
    xt_rsc_0_22_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_22_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_22_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_22_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_22_i_qa_d, xt_rsc_0_22_i_qa_d_bfwt,
      xt_rsc_0_22_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_22_i_bcwt <= '0';
      ELSE
        xt_rsc_0_22_i_bcwt <= NOT((NOT(xt_rsc_0_22_i_bcwt OR xt_rsc_0_22_i_biwt))
            OR xt_rsc_0_22_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_22_i_biwt = '1' ) THEN
        xt_rsc_0_22_i_qa_d_bfwt <= xt_rsc_0_22_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_22_i_oswt : IN STD_LOGIC;
    xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_22_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_22_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_22_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_22_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_22_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_22_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_22_i_bdwt <= xt_rsc_0_22_i_oswt AND core_wen;
  xt_rsc_0_22_i_biwt <= (NOT core_wten) AND xt_rsc_0_22_i_oswt;
  xt_rsc_0_22_i_wea_d_core_sct_pff <= xt_rsc_0_22_i_wea_d_core_psct_pff AND xt_rsc_0_22_i_dswt_pff;
  xt_rsc_0_22_i_dswt_pff <= core_wen AND xt_rsc_0_22_i_oswt_pff;
  xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_22_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_21_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_21_i_biwt : IN STD_LOGIC;
    xt_rsc_0_21_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_21_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_21_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_21_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_21_i_qa_d, xt_rsc_0_21_i_qa_d_bfwt,
      xt_rsc_0_21_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_21_i_bcwt <= '0';
      ELSE
        xt_rsc_0_21_i_bcwt <= NOT((NOT(xt_rsc_0_21_i_bcwt OR xt_rsc_0_21_i_biwt))
            OR xt_rsc_0_21_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_21_i_biwt = '1' ) THEN
        xt_rsc_0_21_i_qa_d_bfwt <= xt_rsc_0_21_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_21_i_oswt : IN STD_LOGIC;
    xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_21_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_21_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_21_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_21_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_21_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_21_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_21_i_bdwt <= xt_rsc_0_21_i_oswt AND core_wen;
  xt_rsc_0_21_i_biwt <= (NOT core_wten) AND xt_rsc_0_21_i_oswt;
  xt_rsc_0_21_i_wea_d_core_sct_pff <= xt_rsc_0_21_i_wea_d_core_psct_pff AND xt_rsc_0_21_i_dswt_pff;
  xt_rsc_0_21_i_dswt_pff <= core_wen AND xt_rsc_0_21_i_oswt_pff;
  xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_21_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_20_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_20_i_biwt : IN STD_LOGIC;
    xt_rsc_0_20_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_20_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_20_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_20_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_20_i_qa_d, xt_rsc_0_20_i_qa_d_bfwt,
      xt_rsc_0_20_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_20_i_bcwt <= '0';
      ELSE
        xt_rsc_0_20_i_bcwt <= NOT((NOT(xt_rsc_0_20_i_bcwt OR xt_rsc_0_20_i_biwt))
            OR xt_rsc_0_20_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_20_i_biwt = '1' ) THEN
        xt_rsc_0_20_i_qa_d_bfwt <= xt_rsc_0_20_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_20_i_oswt : IN STD_LOGIC;
    xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_20_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_20_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_20_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_20_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_20_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_20_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_20_i_bdwt <= xt_rsc_0_20_i_oswt AND core_wen;
  xt_rsc_0_20_i_biwt <= (NOT core_wten) AND xt_rsc_0_20_i_oswt;
  xt_rsc_0_20_i_wea_d_core_sct_pff <= xt_rsc_0_20_i_wea_d_core_psct_pff AND xt_rsc_0_20_i_dswt_pff;
  xt_rsc_0_20_i_dswt_pff <= core_wen AND xt_rsc_0_20_i_oswt_pff;
  xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_20_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_19_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_19_i_biwt : IN STD_LOGIC;
    xt_rsc_0_19_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_19_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_19_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_19_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_19_i_qa_d, xt_rsc_0_19_i_qa_d_bfwt,
      xt_rsc_0_19_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_19_i_bcwt <= '0';
      ELSE
        xt_rsc_0_19_i_bcwt <= NOT((NOT(xt_rsc_0_19_i_bcwt OR xt_rsc_0_19_i_biwt))
            OR xt_rsc_0_19_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_19_i_biwt = '1' ) THEN
        xt_rsc_0_19_i_qa_d_bfwt <= xt_rsc_0_19_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_19_i_oswt : IN STD_LOGIC;
    xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_19_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_19_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_19_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_19_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_19_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_19_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_19_i_bdwt <= xt_rsc_0_19_i_oswt AND core_wen;
  xt_rsc_0_19_i_biwt <= (NOT core_wten) AND xt_rsc_0_19_i_oswt;
  xt_rsc_0_19_i_wea_d_core_sct_pff <= xt_rsc_0_19_i_wea_d_core_psct_pff AND xt_rsc_0_19_i_dswt_pff;
  xt_rsc_0_19_i_dswt_pff <= core_wen AND xt_rsc_0_19_i_oswt_pff;
  xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_19_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_18_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_18_i_biwt : IN STD_LOGIC;
    xt_rsc_0_18_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_18_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_18_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_18_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_18_i_qa_d, xt_rsc_0_18_i_qa_d_bfwt,
      xt_rsc_0_18_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_18_i_bcwt <= '0';
      ELSE
        xt_rsc_0_18_i_bcwt <= NOT((NOT(xt_rsc_0_18_i_bcwt OR xt_rsc_0_18_i_biwt))
            OR xt_rsc_0_18_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_18_i_biwt = '1' ) THEN
        xt_rsc_0_18_i_qa_d_bfwt <= xt_rsc_0_18_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_18_i_oswt : IN STD_LOGIC;
    xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_18_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_18_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_18_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_18_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_18_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_18_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_18_i_bdwt <= xt_rsc_0_18_i_oswt AND core_wen;
  xt_rsc_0_18_i_biwt <= (NOT core_wten) AND xt_rsc_0_18_i_oswt;
  xt_rsc_0_18_i_wea_d_core_sct_pff <= xt_rsc_0_18_i_wea_d_core_psct_pff AND xt_rsc_0_18_i_dswt_pff;
  xt_rsc_0_18_i_dswt_pff <= core_wen AND xt_rsc_0_18_i_oswt_pff;
  xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_18_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_17_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_17_i_biwt : IN STD_LOGIC;
    xt_rsc_0_17_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_17_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_17_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_17_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_17_i_qa_d, xt_rsc_0_17_i_qa_d_bfwt,
      xt_rsc_0_17_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_17_i_bcwt <= '0';
      ELSE
        xt_rsc_0_17_i_bcwt <= NOT((NOT(xt_rsc_0_17_i_bcwt OR xt_rsc_0_17_i_biwt))
            OR xt_rsc_0_17_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_17_i_biwt = '1' ) THEN
        xt_rsc_0_17_i_qa_d_bfwt <= xt_rsc_0_17_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_17_i_oswt : IN STD_LOGIC;
    xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_17_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_17_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_17_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_17_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_17_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_17_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_17_i_bdwt <= xt_rsc_0_17_i_oswt AND core_wen;
  xt_rsc_0_17_i_biwt <= (NOT core_wten) AND xt_rsc_0_17_i_oswt;
  xt_rsc_0_17_i_wea_d_core_sct_pff <= xt_rsc_0_17_i_wea_d_core_psct_pff AND xt_rsc_0_17_i_dswt_pff;
  xt_rsc_0_17_i_dswt_pff <= core_wen AND xt_rsc_0_17_i_oswt_pff;
  xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_17_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_16_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_16_i_biwt : IN STD_LOGIC;
    xt_rsc_0_16_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_16_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_16_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_16_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_16_i_qa_d, xt_rsc_0_16_i_qa_d_bfwt,
      xt_rsc_0_16_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_16_i_bcwt <= '0';
      ELSE
        xt_rsc_0_16_i_bcwt <= NOT((NOT(xt_rsc_0_16_i_bcwt OR xt_rsc_0_16_i_biwt))
            OR xt_rsc_0_16_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_16_i_biwt = '1' ) THEN
        xt_rsc_0_16_i_qa_d_bfwt <= xt_rsc_0_16_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_16_i_oswt : IN STD_LOGIC;
    xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_16_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_16_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_16_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_16_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_16_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_16_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_16_i_bdwt <= xt_rsc_0_16_i_oswt AND core_wen;
  xt_rsc_0_16_i_biwt <= (NOT core_wten) AND xt_rsc_0_16_i_oswt;
  xt_rsc_0_16_i_wea_d_core_sct_pff <= xt_rsc_0_16_i_wea_d_core_psct_pff AND xt_rsc_0_16_i_dswt_pff;
  xt_rsc_0_16_i_dswt_pff <= core_wen AND xt_rsc_0_16_i_oswt_pff;
  xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_16_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_15_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_15_i_biwt : IN STD_LOGIC;
    xt_rsc_0_15_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_15_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_15_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_15_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_15_i_qa_d, xt_rsc_0_15_i_qa_d_bfwt,
      xt_rsc_0_15_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_15_i_bcwt <= '0';
      ELSE
        xt_rsc_0_15_i_bcwt <= NOT((NOT(xt_rsc_0_15_i_bcwt OR xt_rsc_0_15_i_biwt))
            OR xt_rsc_0_15_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_15_i_biwt = '1' ) THEN
        xt_rsc_0_15_i_qa_d_bfwt <= xt_rsc_0_15_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_15_i_oswt : IN STD_LOGIC;
    xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_15_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_15_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_15_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_15_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_15_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_15_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_15_i_bdwt <= xt_rsc_0_15_i_oswt AND core_wen;
  xt_rsc_0_15_i_biwt <= (NOT core_wten) AND xt_rsc_0_15_i_oswt;
  xt_rsc_0_15_i_wea_d_core_sct_pff <= xt_rsc_0_15_i_wea_d_core_psct_pff AND xt_rsc_0_15_i_dswt_pff;
  xt_rsc_0_15_i_dswt_pff <= core_wen AND xt_rsc_0_15_i_oswt_pff;
  xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_15_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_14_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_14_i_biwt : IN STD_LOGIC;
    xt_rsc_0_14_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_14_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_14_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_14_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_14_i_qa_d, xt_rsc_0_14_i_qa_d_bfwt,
      xt_rsc_0_14_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_14_i_bcwt <= '0';
      ELSE
        xt_rsc_0_14_i_bcwt <= NOT((NOT(xt_rsc_0_14_i_bcwt OR xt_rsc_0_14_i_biwt))
            OR xt_rsc_0_14_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_14_i_biwt = '1' ) THEN
        xt_rsc_0_14_i_qa_d_bfwt <= xt_rsc_0_14_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_14_i_oswt : IN STD_LOGIC;
    xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_14_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_14_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_14_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_14_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_14_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_14_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_14_i_bdwt <= xt_rsc_0_14_i_oswt AND core_wen;
  xt_rsc_0_14_i_biwt <= (NOT core_wten) AND xt_rsc_0_14_i_oswt;
  xt_rsc_0_14_i_wea_d_core_sct_pff <= xt_rsc_0_14_i_wea_d_core_psct_pff AND xt_rsc_0_14_i_dswt_pff;
  xt_rsc_0_14_i_dswt_pff <= core_wen AND xt_rsc_0_14_i_oswt_pff;
  xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_14_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_13_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_13_i_biwt : IN STD_LOGIC;
    xt_rsc_0_13_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_13_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_13_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_13_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_13_i_qa_d, xt_rsc_0_13_i_qa_d_bfwt,
      xt_rsc_0_13_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_13_i_bcwt <= '0';
      ELSE
        xt_rsc_0_13_i_bcwt <= NOT((NOT(xt_rsc_0_13_i_bcwt OR xt_rsc_0_13_i_biwt))
            OR xt_rsc_0_13_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_13_i_biwt = '1' ) THEN
        xt_rsc_0_13_i_qa_d_bfwt <= xt_rsc_0_13_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_13_i_oswt : IN STD_LOGIC;
    xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_13_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_13_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_13_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_13_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_13_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_13_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_13_i_bdwt <= xt_rsc_0_13_i_oswt AND core_wen;
  xt_rsc_0_13_i_biwt <= (NOT core_wten) AND xt_rsc_0_13_i_oswt;
  xt_rsc_0_13_i_wea_d_core_sct_pff <= xt_rsc_0_13_i_wea_d_core_psct_pff AND xt_rsc_0_13_i_dswt_pff;
  xt_rsc_0_13_i_dswt_pff <= core_wen AND xt_rsc_0_13_i_oswt_pff;
  xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_13_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_12_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_12_i_biwt : IN STD_LOGIC;
    xt_rsc_0_12_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_12_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_12_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_12_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_12_i_qa_d, xt_rsc_0_12_i_qa_d_bfwt,
      xt_rsc_0_12_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_12_i_bcwt <= '0';
      ELSE
        xt_rsc_0_12_i_bcwt <= NOT((NOT(xt_rsc_0_12_i_bcwt OR xt_rsc_0_12_i_biwt))
            OR xt_rsc_0_12_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_12_i_biwt = '1' ) THEN
        xt_rsc_0_12_i_qa_d_bfwt <= xt_rsc_0_12_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_12_i_oswt : IN STD_LOGIC;
    xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_12_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_12_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_12_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_12_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_12_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_12_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_12_i_bdwt <= xt_rsc_0_12_i_oswt AND core_wen;
  xt_rsc_0_12_i_biwt <= (NOT core_wten) AND xt_rsc_0_12_i_oswt;
  xt_rsc_0_12_i_wea_d_core_sct_pff <= xt_rsc_0_12_i_wea_d_core_psct_pff AND xt_rsc_0_12_i_dswt_pff;
  xt_rsc_0_12_i_dswt_pff <= core_wen AND xt_rsc_0_12_i_oswt_pff;
  xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_12_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_11_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_11_i_biwt : IN STD_LOGIC;
    xt_rsc_0_11_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_11_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_11_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_11_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_11_i_qa_d, xt_rsc_0_11_i_qa_d_bfwt,
      xt_rsc_0_11_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_11_i_bcwt <= '0';
      ELSE
        xt_rsc_0_11_i_bcwt <= NOT((NOT(xt_rsc_0_11_i_bcwt OR xt_rsc_0_11_i_biwt))
            OR xt_rsc_0_11_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_11_i_biwt = '1' ) THEN
        xt_rsc_0_11_i_qa_d_bfwt <= xt_rsc_0_11_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_11_i_oswt : IN STD_LOGIC;
    xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_11_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_11_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_11_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_11_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_11_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_11_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_11_i_bdwt <= xt_rsc_0_11_i_oswt AND core_wen;
  xt_rsc_0_11_i_biwt <= (NOT core_wten) AND xt_rsc_0_11_i_oswt;
  xt_rsc_0_11_i_wea_d_core_sct_pff <= xt_rsc_0_11_i_wea_d_core_psct_pff AND xt_rsc_0_11_i_dswt_pff;
  xt_rsc_0_11_i_dswt_pff <= core_wen AND xt_rsc_0_11_i_oswt_pff;
  xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_11_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_10_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_10_i_biwt : IN STD_LOGIC;
    xt_rsc_0_10_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_10_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_10_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_10_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_10_i_qa_d, xt_rsc_0_10_i_qa_d_bfwt,
      xt_rsc_0_10_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_10_i_bcwt <= '0';
      ELSE
        xt_rsc_0_10_i_bcwt <= NOT((NOT(xt_rsc_0_10_i_bcwt OR xt_rsc_0_10_i_biwt))
            OR xt_rsc_0_10_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_10_i_biwt = '1' ) THEN
        xt_rsc_0_10_i_qa_d_bfwt <= xt_rsc_0_10_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_10_i_oswt : IN STD_LOGIC;
    xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_10_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_10_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_10_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_10_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_10_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_10_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_10_i_bdwt <= xt_rsc_0_10_i_oswt AND core_wen;
  xt_rsc_0_10_i_biwt <= (NOT core_wten) AND xt_rsc_0_10_i_oswt;
  xt_rsc_0_10_i_wea_d_core_sct_pff <= xt_rsc_0_10_i_wea_d_core_psct_pff AND xt_rsc_0_10_i_dswt_pff;
  xt_rsc_0_10_i_dswt_pff <= core_wen AND xt_rsc_0_10_i_oswt_pff;
  xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_10_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_9_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_9_i_biwt : IN STD_LOGIC;
    xt_rsc_0_9_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_9_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_9_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_9_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_9_i_qa_d, xt_rsc_0_9_i_qa_d_bfwt,
      xt_rsc_0_9_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_9_i_bcwt <= '0';
      ELSE
        xt_rsc_0_9_i_bcwt <= NOT((NOT(xt_rsc_0_9_i_bcwt OR xt_rsc_0_9_i_biwt)) OR
            xt_rsc_0_9_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_9_i_biwt = '1' ) THEN
        xt_rsc_0_9_i_qa_d_bfwt <= xt_rsc_0_9_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_9_i_oswt : IN STD_LOGIC;
    xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_9_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_9_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_9_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_9_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_9_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_9_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_9_i_bdwt <= xt_rsc_0_9_i_oswt AND core_wen;
  xt_rsc_0_9_i_biwt <= (NOT core_wten) AND xt_rsc_0_9_i_oswt;
  xt_rsc_0_9_i_wea_d_core_sct_pff <= xt_rsc_0_9_i_wea_d_core_psct_pff AND xt_rsc_0_9_i_dswt_pff;
  xt_rsc_0_9_i_dswt_pff <= core_wen AND xt_rsc_0_9_i_oswt_pff;
  xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_9_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_8_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_8_i_biwt : IN STD_LOGIC;
    xt_rsc_0_8_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_8_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_8_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_8_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_8_i_qa_d, xt_rsc_0_8_i_qa_d_bfwt,
      xt_rsc_0_8_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_8_i_bcwt <= '0';
      ELSE
        xt_rsc_0_8_i_bcwt <= NOT((NOT(xt_rsc_0_8_i_bcwt OR xt_rsc_0_8_i_biwt)) OR
            xt_rsc_0_8_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_8_i_biwt = '1' ) THEN
        xt_rsc_0_8_i_qa_d_bfwt <= xt_rsc_0_8_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_8_i_oswt : IN STD_LOGIC;
    xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_8_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_8_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_8_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_8_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_8_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_8_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_8_i_bdwt <= xt_rsc_0_8_i_oswt AND core_wen;
  xt_rsc_0_8_i_biwt <= (NOT core_wten) AND xt_rsc_0_8_i_oswt;
  xt_rsc_0_8_i_wea_d_core_sct_pff <= xt_rsc_0_8_i_wea_d_core_psct_pff AND xt_rsc_0_8_i_dswt_pff;
  xt_rsc_0_8_i_dswt_pff <= core_wen AND xt_rsc_0_8_i_oswt_pff;
  xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_8_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_7_i_biwt : IN STD_LOGIC;
    xt_rsc_0_7_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_7_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_7_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_7_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_7_i_qa_d, xt_rsc_0_7_i_qa_d_bfwt,
      xt_rsc_0_7_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_7_i_bcwt <= '0';
      ELSE
        xt_rsc_0_7_i_bcwt <= NOT((NOT(xt_rsc_0_7_i_bcwt OR xt_rsc_0_7_i_biwt)) OR
            xt_rsc_0_7_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_7_i_biwt = '1' ) THEN
        xt_rsc_0_7_i_qa_d_bfwt <= xt_rsc_0_7_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_7_i_oswt : IN STD_LOGIC;
    xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_7_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_7_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_7_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_7_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_7_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_7_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_7_i_bdwt <= xt_rsc_0_7_i_oswt AND core_wen;
  xt_rsc_0_7_i_biwt <= (NOT core_wten) AND xt_rsc_0_7_i_oswt;
  xt_rsc_0_7_i_wea_d_core_sct_pff <= xt_rsc_0_7_i_wea_d_core_psct_pff AND xt_rsc_0_7_i_dswt_pff;
  xt_rsc_0_7_i_dswt_pff <= core_wen AND xt_rsc_0_7_i_oswt_pff;
  xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_7_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_6_i_biwt : IN STD_LOGIC;
    xt_rsc_0_6_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_6_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_6_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_6_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_6_i_qa_d, xt_rsc_0_6_i_qa_d_bfwt,
      xt_rsc_0_6_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_6_i_bcwt <= '0';
      ELSE
        xt_rsc_0_6_i_bcwt <= NOT((NOT(xt_rsc_0_6_i_bcwt OR xt_rsc_0_6_i_biwt)) OR
            xt_rsc_0_6_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_6_i_biwt = '1' ) THEN
        xt_rsc_0_6_i_qa_d_bfwt <= xt_rsc_0_6_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_6_i_oswt : IN STD_LOGIC;
    xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_6_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_6_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_6_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_6_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_6_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_6_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_6_i_bdwt <= xt_rsc_0_6_i_oswt AND core_wen;
  xt_rsc_0_6_i_biwt <= (NOT core_wten) AND xt_rsc_0_6_i_oswt;
  xt_rsc_0_6_i_wea_d_core_sct_pff <= xt_rsc_0_6_i_wea_d_core_psct_pff AND xt_rsc_0_6_i_dswt_pff;
  xt_rsc_0_6_i_dswt_pff <= core_wen AND xt_rsc_0_6_i_oswt_pff;
  xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_6_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_5_i_biwt : IN STD_LOGIC;
    xt_rsc_0_5_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_5_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_5_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_5_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_5_i_qa_d, xt_rsc_0_5_i_qa_d_bfwt,
      xt_rsc_0_5_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_5_i_bcwt <= '0';
      ELSE
        xt_rsc_0_5_i_bcwt <= NOT((NOT(xt_rsc_0_5_i_bcwt OR xt_rsc_0_5_i_biwt)) OR
            xt_rsc_0_5_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_5_i_biwt = '1' ) THEN
        xt_rsc_0_5_i_qa_d_bfwt <= xt_rsc_0_5_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_5_i_oswt : IN STD_LOGIC;
    xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_5_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_5_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_5_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_5_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_5_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_5_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_5_i_bdwt <= xt_rsc_0_5_i_oswt AND core_wen;
  xt_rsc_0_5_i_biwt <= (NOT core_wten) AND xt_rsc_0_5_i_oswt;
  xt_rsc_0_5_i_wea_d_core_sct_pff <= xt_rsc_0_5_i_wea_d_core_psct_pff AND xt_rsc_0_5_i_dswt_pff;
  xt_rsc_0_5_i_dswt_pff <= core_wen AND xt_rsc_0_5_i_oswt_pff;
  xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_5_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_4_i_biwt : IN STD_LOGIC;
    xt_rsc_0_4_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_4_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_4_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_4_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_4_i_qa_d, xt_rsc_0_4_i_qa_d_bfwt,
      xt_rsc_0_4_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_4_i_bcwt <= '0';
      ELSE
        xt_rsc_0_4_i_bcwt <= NOT((NOT(xt_rsc_0_4_i_bcwt OR xt_rsc_0_4_i_biwt)) OR
            xt_rsc_0_4_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_4_i_biwt = '1' ) THEN
        xt_rsc_0_4_i_qa_d_bfwt <= xt_rsc_0_4_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_4_i_oswt : IN STD_LOGIC;
    xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_4_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_4_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_4_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_4_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_4_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_4_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_4_i_bdwt <= xt_rsc_0_4_i_oswt AND core_wen;
  xt_rsc_0_4_i_biwt <= (NOT core_wten) AND xt_rsc_0_4_i_oswt;
  xt_rsc_0_4_i_wea_d_core_sct_pff <= xt_rsc_0_4_i_wea_d_core_psct_pff AND xt_rsc_0_4_i_dswt_pff;
  xt_rsc_0_4_i_dswt_pff <= core_wen AND xt_rsc_0_4_i_oswt_pff;
  xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_4_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_3_i_biwt : IN STD_LOGIC;
    xt_rsc_0_3_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_3_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_3_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_3_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_3_i_qa_d, xt_rsc_0_3_i_qa_d_bfwt,
      xt_rsc_0_3_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_3_i_bcwt <= '0';
      ELSE
        xt_rsc_0_3_i_bcwt <= NOT((NOT(xt_rsc_0_3_i_bcwt OR xt_rsc_0_3_i_biwt)) OR
            xt_rsc_0_3_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_3_i_biwt = '1' ) THEN
        xt_rsc_0_3_i_qa_d_bfwt <= xt_rsc_0_3_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_3_i_oswt : IN STD_LOGIC;
    xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_3_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_3_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_3_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_3_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_3_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_3_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_3_i_bdwt <= xt_rsc_0_3_i_oswt AND core_wen;
  xt_rsc_0_3_i_biwt <= (NOT core_wten) AND xt_rsc_0_3_i_oswt;
  xt_rsc_0_3_i_wea_d_core_sct_pff <= xt_rsc_0_3_i_wea_d_core_psct_pff AND xt_rsc_0_3_i_dswt_pff;
  xt_rsc_0_3_i_dswt_pff <= core_wen AND xt_rsc_0_3_i_oswt_pff;
  xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_3_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_2_i_biwt : IN STD_LOGIC;
    xt_rsc_0_2_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_2_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_2_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_2_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_2_i_qa_d, xt_rsc_0_2_i_qa_d_bfwt,
      xt_rsc_0_2_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_2_i_bcwt <= '0';
      ELSE
        xt_rsc_0_2_i_bcwt <= NOT((NOT(xt_rsc_0_2_i_bcwt OR xt_rsc_0_2_i_biwt)) OR
            xt_rsc_0_2_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_2_i_biwt = '1' ) THEN
        xt_rsc_0_2_i_qa_d_bfwt <= xt_rsc_0_2_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_2_i_oswt : IN STD_LOGIC;
    xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_2_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_2_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_2_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_2_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_2_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_2_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_2_i_bdwt <= xt_rsc_0_2_i_oswt AND core_wen;
  xt_rsc_0_2_i_biwt <= (NOT core_wten) AND xt_rsc_0_2_i_oswt;
  xt_rsc_0_2_i_wea_d_core_sct_pff <= xt_rsc_0_2_i_wea_d_core_psct_pff AND xt_rsc_0_2_i_dswt_pff;
  xt_rsc_0_2_i_dswt_pff <= core_wen AND xt_rsc_0_2_i_oswt_pff;
  xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_2_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_1_i_biwt : IN STD_LOGIC;
    xt_rsc_0_1_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_1_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_1_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_1_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_1_i_qa_d, xt_rsc_0_1_i_qa_d_bfwt,
      xt_rsc_0_1_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_1_i_bcwt <= '0';
      ELSE
        xt_rsc_0_1_i_bcwt <= NOT((NOT(xt_rsc_0_1_i_bcwt OR xt_rsc_0_1_i_biwt)) OR
            xt_rsc_0_1_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_1_i_biwt = '1' ) THEN
        xt_rsc_0_1_i_qa_d_bfwt <= xt_rsc_0_1_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_1_i_oswt : IN STD_LOGIC;
    xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_1_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_1_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_1_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_1_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_1_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_1_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_1_i_bdwt <= xt_rsc_0_1_i_oswt AND core_wen;
  xt_rsc_0_1_i_biwt <= (NOT core_wten) AND xt_rsc_0_1_i_oswt;
  xt_rsc_0_1_i_wea_d_core_sct_pff <= xt_rsc_0_1_i_wea_d_core_psct_pff AND xt_rsc_0_1_i_dswt_pff;
  xt_rsc_0_1_i_dswt_pff <= core_wen AND xt_rsc_0_1_i_oswt_pff;
  xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_1_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_dp IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_0_i_biwt : IN STD_LOGIC;
    xt_rsc_0_0_i_bdwt : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_dp IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_0_i_bcwt : STD_LOGIC;
  SIGNAL xt_rsc_0_0_i_qa_d_bfwt : STD_LOGIC_VECTOR (31 DOWNTO 0);

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  xt_rsc_0_0_i_qa_d_mxwt <= MUX_v_32_2_2(xt_rsc_0_0_i_qa_d, xt_rsc_0_0_i_qa_d_bfwt,
      xt_rsc_0_0_i_bcwt);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        xt_rsc_0_0_i_bcwt <= '0';
      ELSE
        xt_rsc_0_0_i_bcwt <= NOT((NOT(xt_rsc_0_0_i_bcwt OR xt_rsc_0_0_i_biwt)) OR
            xt_rsc_0_0_i_bdwt);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( xt_rsc_0_0_i_biwt = '1' ) THEN
        xt_rsc_0_0_i_qa_d_bfwt <= xt_rsc_0_0_i_qa_d;
      END IF;
    END IF;
  END PROCESS;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_ctrl
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_ctrl IS
  PORT(
    core_wen : IN STD_LOGIC;
    xt_rsc_0_0_i_oswt : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_0_i_biwt : OUT STD_LOGIC;
    xt_rsc_0_0_i_bdwt : OUT STD_LOGIC;
    xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
    xt_rsc_0_0_i_wea_d_core_sct_pff : OUT STD_LOGIC;
    xt_rsc_0_0_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_0_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_ctrl;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_ctrl IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_0_i_dswt_pff : STD_LOGIC;

BEGIN
  xt_rsc_0_0_i_bdwt <= xt_rsc_0_0_i_oswt AND core_wen;
  xt_rsc_0_0_i_biwt <= (NOT core_wten) AND xt_rsc_0_0_i_oswt;
  xt_rsc_0_0_i_wea_d_core_sct_pff <= xt_rsc_0_0_i_wea_d_core_psct_pff AND xt_rsc_0_0_i_dswt_pff;
  xt_rsc_0_0_i_dswt_pff <= core_wen AND xt_rsc_0_0_i_oswt_pff;
  xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct <= xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct
      AND xt_rsc_0_0_i_dswt_pff;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_wait_dp
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_wait_dp IS
  PORT(
    yt_rsc_0_0_cgo_iro : IN STD_LOGIC;
    yt_rsc_0_0_i_clken_d : OUT STD_LOGIC;
    yt_rsc_0_16_cgo_iro : IN STD_LOGIC;
    yt_rsc_0_16_i_clken_d : OUT STD_LOGIC;
    yt_rsc_1_0_cgo_iro : IN STD_LOGIC;
    yt_rsc_1_0_i_clken_d : OUT STD_LOGIC;
    yt_rsc_1_16_cgo_iro : IN STD_LOGIC;
    yt_rsc_1_16_i_clken_d : OUT STD_LOGIC;
    ensig_cgo_iro : IN STD_LOGIC;
    ensig_cgo_iro_17 : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    yt_rsc_0_0_cgo : IN STD_LOGIC;
    yt_rsc_0_16_cgo : IN STD_LOGIC;
    yt_rsc_1_0_cgo : IN STD_LOGIC;
    yt_rsc_1_16_cgo : IN STD_LOGIC;
    ensig_cgo : IN STD_LOGIC;
    mult_t_mul_cmp_en : OUT STD_LOGIC;
    ensig_cgo_17 : IN STD_LOGIC;
    mult_z_mul_cmp_1_en : OUT STD_LOGIC
  );
END peaseNTT_core_wait_dp;

ARCHITECTURE v29 OF peaseNTT_core_wait_dp IS
  -- Default Constants

BEGIN
  yt_rsc_0_0_i_clken_d <= core_wen AND (yt_rsc_0_0_cgo OR yt_rsc_0_0_cgo_iro);
  yt_rsc_0_16_i_clken_d <= core_wen AND (yt_rsc_0_16_cgo OR yt_rsc_0_16_cgo_iro);
  yt_rsc_1_0_i_clken_d <= core_wen AND (yt_rsc_1_0_cgo OR yt_rsc_1_0_cgo_iro);
  yt_rsc_1_16_i_clken_d <= core_wen AND (yt_rsc_1_16_cgo OR yt_rsc_1_16_cgo_iro);
  mult_t_mul_cmp_en <= core_wen AND (ensig_cgo OR ensig_cgo_iro);
  mult_z_mul_cmp_1_en <= core_wen AND (ensig_cgo_17 OR ensig_cgo_iro_17);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_0_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_0_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_0_obj_twiddle_h_rsc_triosy_0_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_0_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_0_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_0_obj_twiddle_h_rsc_triosy_0_0_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_0_obj_twiddle_h_rsc_triosy_0_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_0_obj_iswt0 => twiddle_h_rsc_triosy_0_0_obj_iswt0,
      twiddle_h_rsc_triosy_0_0_obj_ld_core_sct => twiddle_h_rsc_triosy_0_0_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_1_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_1_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_1_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_1_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_1_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_1_obj_twiddle_h_rsc_triosy_0_1_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_1_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_1_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_1_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_1_obj_twiddle_h_rsc_triosy_0_1_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_1_obj_twiddle_h_rsc_triosy_0_1_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_1_obj_iswt0 => twiddle_h_rsc_triosy_0_1_obj_iswt0,
      twiddle_h_rsc_triosy_0_1_obj_ld_core_sct => twiddle_h_rsc_triosy_0_1_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_2_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_2_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_2_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_2_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_2_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_2_obj_twiddle_h_rsc_triosy_0_2_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_2_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_2_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_2_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_2_obj_twiddle_h_rsc_triosy_0_2_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_2_obj_twiddle_h_rsc_triosy_0_2_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_2_obj_iswt0 => twiddle_h_rsc_triosy_0_2_obj_iswt0,
      twiddle_h_rsc_triosy_0_2_obj_ld_core_sct => twiddle_h_rsc_triosy_0_2_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_3_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_3_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_3_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_3_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_3_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_3_obj_twiddle_h_rsc_triosy_0_3_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_3_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_3_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_3_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_3_obj_twiddle_h_rsc_triosy_0_3_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_3_obj_twiddle_h_rsc_triosy_0_3_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_3_obj_iswt0 => twiddle_h_rsc_triosy_0_3_obj_iswt0,
      twiddle_h_rsc_triosy_0_3_obj_ld_core_sct => twiddle_h_rsc_triosy_0_3_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_4_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_4_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_4_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_4_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_4_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_4_obj_twiddle_h_rsc_triosy_0_4_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_4_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_4_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_4_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_4_obj_twiddle_h_rsc_triosy_0_4_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_4_obj_twiddle_h_rsc_triosy_0_4_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_4_obj_iswt0 => twiddle_h_rsc_triosy_0_4_obj_iswt0,
      twiddle_h_rsc_triosy_0_4_obj_ld_core_sct => twiddle_h_rsc_triosy_0_4_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_5_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_5_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_5_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_5_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_5_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_5_obj_twiddle_h_rsc_triosy_0_5_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_5_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_5_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_5_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_5_obj_twiddle_h_rsc_triosy_0_5_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_5_obj_twiddle_h_rsc_triosy_0_5_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_5_obj_iswt0 => twiddle_h_rsc_triosy_0_5_obj_iswt0,
      twiddle_h_rsc_triosy_0_5_obj_ld_core_sct => twiddle_h_rsc_triosy_0_5_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_6_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_6_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_6_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_6_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_6_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_6_obj_twiddle_h_rsc_triosy_0_6_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_6_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_6_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_6_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_6_obj_twiddle_h_rsc_triosy_0_6_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_6_obj_twiddle_h_rsc_triosy_0_6_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_6_obj_iswt0 => twiddle_h_rsc_triosy_0_6_obj_iswt0,
      twiddle_h_rsc_triosy_0_6_obj_ld_core_sct => twiddle_h_rsc_triosy_0_6_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_7_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_7_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_7_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_7_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_7_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_7_obj_twiddle_h_rsc_triosy_0_7_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_7_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_7_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_7_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_7_obj_twiddle_h_rsc_triosy_0_7_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_7_obj_twiddle_h_rsc_triosy_0_7_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_7_obj_iswt0 => twiddle_h_rsc_triosy_0_7_obj_iswt0,
      twiddle_h_rsc_triosy_0_7_obj_ld_core_sct => twiddle_h_rsc_triosy_0_7_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_8_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_8_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_8_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_8_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_8_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_8_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_8_obj_twiddle_h_rsc_triosy_0_8_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_8_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_8_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_8_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_8_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_8_obj_twiddle_h_rsc_triosy_0_8_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_8_obj_twiddle_h_rsc_triosy_0_8_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_8_obj_iswt0 => twiddle_h_rsc_triosy_0_8_obj_iswt0,
      twiddle_h_rsc_triosy_0_8_obj_ld_core_sct => twiddle_h_rsc_triosy_0_8_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_9_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_9_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_9_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_9_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_9_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_9_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_9_obj_twiddle_h_rsc_triosy_0_9_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_9_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_9_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_9_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_9_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_9_obj_twiddle_h_rsc_triosy_0_9_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_9_obj_twiddle_h_rsc_triosy_0_9_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_9_obj_iswt0 => twiddle_h_rsc_triosy_0_9_obj_iswt0,
      twiddle_h_rsc_triosy_0_9_obj_ld_core_sct => twiddle_h_rsc_triosy_0_9_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_10_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_10_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_10_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_10_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_10_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_10_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_10_obj_twiddle_h_rsc_triosy_0_10_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_10_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_10_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_10_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_10_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_10_obj_twiddle_h_rsc_triosy_0_10_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_10_obj_twiddle_h_rsc_triosy_0_10_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_10_obj_iswt0 => twiddle_h_rsc_triosy_0_10_obj_iswt0,
      twiddle_h_rsc_triosy_0_10_obj_ld_core_sct => twiddle_h_rsc_triosy_0_10_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_11_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_11_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_11_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_11_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_11_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_11_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_11_obj_twiddle_h_rsc_triosy_0_11_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_11_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_11_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_11_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_11_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_11_obj_twiddle_h_rsc_triosy_0_11_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_11_obj_twiddle_h_rsc_triosy_0_11_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_11_obj_iswt0 => twiddle_h_rsc_triosy_0_11_obj_iswt0,
      twiddle_h_rsc_triosy_0_11_obj_ld_core_sct => twiddle_h_rsc_triosy_0_11_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_12_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_12_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_12_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_12_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_12_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_12_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_12_obj_twiddle_h_rsc_triosy_0_12_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_12_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_12_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_12_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_12_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_12_obj_twiddle_h_rsc_triosy_0_12_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_12_obj_twiddle_h_rsc_triosy_0_12_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_12_obj_iswt0 => twiddle_h_rsc_triosy_0_12_obj_iswt0,
      twiddle_h_rsc_triosy_0_12_obj_ld_core_sct => twiddle_h_rsc_triosy_0_12_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_13_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_13_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_13_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_13_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_13_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_13_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_13_obj_twiddle_h_rsc_triosy_0_13_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_13_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_13_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_13_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_13_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_13_obj_twiddle_h_rsc_triosy_0_13_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_13_obj_twiddle_h_rsc_triosy_0_13_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_13_obj_iswt0 => twiddle_h_rsc_triosy_0_13_obj_iswt0,
      twiddle_h_rsc_triosy_0_13_obj_ld_core_sct => twiddle_h_rsc_triosy_0_13_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_14_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_14_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_14_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_14_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_14_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_14_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_14_obj_twiddle_h_rsc_triosy_0_14_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_14_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_14_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_14_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_14_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_14_obj_twiddle_h_rsc_triosy_0_14_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_14_obj_twiddle_h_rsc_triosy_0_14_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_14_obj_iswt0 => twiddle_h_rsc_triosy_0_14_obj_iswt0,
      twiddle_h_rsc_triosy_0_14_obj_ld_core_sct => twiddle_h_rsc_triosy_0_14_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_triosy_0_15_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_triosy_0_15_obj IS
  PORT(
    twiddle_h_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_15_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_h_rsc_triosy_0_15_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_triosy_0_15_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_triosy_0_15_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_15_obj_twiddle_h_rsc_triosy_0_15_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_15_obj_iswt0 : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_15_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_h_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_h_rsc_triosy_0_15_obj_ld_core_sct,
      lz => twiddle_h_rsc_triosy_0_15_lz
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_15_obj_twiddle_h_rsc_triosy_0_15_wait_ctrl_inst
      : peaseNTT_core_twiddle_h_rsc_triosy_0_15_obj_twiddle_h_rsc_triosy_0_15_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_15_obj_iswt0 => twiddle_h_rsc_triosy_0_15_obj_iswt0,
      twiddle_h_rsc_triosy_0_15_obj_ld_core_sct => twiddle_h_rsc_triosy_0_15_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_0_obj IS
  PORT(
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_0_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_0_obj_twiddle_rsc_triosy_0_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_0_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_0_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_0_obj_twiddle_rsc_triosy_0_0_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_0_obj_twiddle_rsc_triosy_0_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_0_obj_iswt0 => twiddle_rsc_triosy_0_0_obj_iswt0,
      twiddle_rsc_triosy_0_0_obj_ld_core_sct => twiddle_rsc_triosy_0_0_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_1_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_1_obj IS
  PORT(
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_1_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_1_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_1_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_1_obj_twiddle_rsc_triosy_0_1_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_1_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_1_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_1_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_1_obj_twiddle_rsc_triosy_0_1_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_1_obj_twiddle_rsc_triosy_0_1_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_1_obj_iswt0 => twiddle_rsc_triosy_0_1_obj_iswt0,
      twiddle_rsc_triosy_0_1_obj_ld_core_sct => twiddle_rsc_triosy_0_1_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_2_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_2_obj IS
  PORT(
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_2_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_2_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_2_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_2_obj_twiddle_rsc_triosy_0_2_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_2_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_2_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_2_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_2_obj_twiddle_rsc_triosy_0_2_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_2_obj_twiddle_rsc_triosy_0_2_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_2_obj_iswt0 => twiddle_rsc_triosy_0_2_obj_iswt0,
      twiddle_rsc_triosy_0_2_obj_ld_core_sct => twiddle_rsc_triosy_0_2_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_3_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_3_obj IS
  PORT(
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_3_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_3_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_3_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_3_obj_twiddle_rsc_triosy_0_3_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_3_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_3_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_3_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_3_obj_twiddle_rsc_triosy_0_3_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_3_obj_twiddle_rsc_triosy_0_3_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_3_obj_iswt0 => twiddle_rsc_triosy_0_3_obj_iswt0,
      twiddle_rsc_triosy_0_3_obj_ld_core_sct => twiddle_rsc_triosy_0_3_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_4_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_4_obj IS
  PORT(
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_4_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_4_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_4_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_4_obj_twiddle_rsc_triosy_0_4_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_4_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_4_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_4_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_4_obj_twiddle_rsc_triosy_0_4_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_4_obj_twiddle_rsc_triosy_0_4_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_4_obj_iswt0 => twiddle_rsc_triosy_0_4_obj_iswt0,
      twiddle_rsc_triosy_0_4_obj_ld_core_sct => twiddle_rsc_triosy_0_4_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_5_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_5_obj IS
  PORT(
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_5_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_5_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_5_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_5_obj_twiddle_rsc_triosy_0_5_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_5_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_5_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_5_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_5_obj_twiddle_rsc_triosy_0_5_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_5_obj_twiddle_rsc_triosy_0_5_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_5_obj_iswt0 => twiddle_rsc_triosy_0_5_obj_iswt0,
      twiddle_rsc_triosy_0_5_obj_ld_core_sct => twiddle_rsc_triosy_0_5_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_6_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_6_obj IS
  PORT(
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_6_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_6_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_6_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_6_obj_twiddle_rsc_triosy_0_6_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_6_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_6_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_6_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_6_obj_twiddle_rsc_triosy_0_6_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_6_obj_twiddle_rsc_triosy_0_6_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_6_obj_iswt0 => twiddle_rsc_triosy_0_6_obj_iswt0,
      twiddle_rsc_triosy_0_6_obj_ld_core_sct => twiddle_rsc_triosy_0_6_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_7_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_7_obj IS
  PORT(
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_7_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_7_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_7_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_7_obj_twiddle_rsc_triosy_0_7_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_7_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_7_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_7_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_7_obj_twiddle_rsc_triosy_0_7_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_7_obj_twiddle_rsc_triosy_0_7_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_7_obj_iswt0 => twiddle_rsc_triosy_0_7_obj_iswt0,
      twiddle_rsc_triosy_0_7_obj_ld_core_sct => twiddle_rsc_triosy_0_7_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_8_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_8_obj IS
  PORT(
    twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_8_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_8_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_8_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_8_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_8_obj_twiddle_rsc_triosy_0_8_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_8_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_8_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_8_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_8_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_8_obj_twiddle_rsc_triosy_0_8_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_8_obj_twiddle_rsc_triosy_0_8_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_8_obj_iswt0 => twiddle_rsc_triosy_0_8_obj_iswt0,
      twiddle_rsc_triosy_0_8_obj_ld_core_sct => twiddle_rsc_triosy_0_8_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_9_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_9_obj IS
  PORT(
    twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_9_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_9_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_9_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_9_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_9_obj_twiddle_rsc_triosy_0_9_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_9_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_9_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_9_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_9_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_9_obj_twiddle_rsc_triosy_0_9_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_9_obj_twiddle_rsc_triosy_0_9_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_9_obj_iswt0 => twiddle_rsc_triosy_0_9_obj_iswt0,
      twiddle_rsc_triosy_0_9_obj_ld_core_sct => twiddle_rsc_triosy_0_9_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_10_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_10_obj IS
  PORT(
    twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_10_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_10_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_10_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_10_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_10_obj_twiddle_rsc_triosy_0_10_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_10_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_10_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_10_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_10_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_10_obj_twiddle_rsc_triosy_0_10_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_10_obj_twiddle_rsc_triosy_0_10_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_10_obj_iswt0 => twiddle_rsc_triosy_0_10_obj_iswt0,
      twiddle_rsc_triosy_0_10_obj_ld_core_sct => twiddle_rsc_triosy_0_10_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_11_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_11_obj IS
  PORT(
    twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_11_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_11_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_11_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_11_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_11_obj_twiddle_rsc_triosy_0_11_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_11_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_11_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_11_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_11_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_11_obj_twiddle_rsc_triosy_0_11_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_11_obj_twiddle_rsc_triosy_0_11_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_11_obj_iswt0 => twiddle_rsc_triosy_0_11_obj_iswt0,
      twiddle_rsc_triosy_0_11_obj_ld_core_sct => twiddle_rsc_triosy_0_11_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_12_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_12_obj IS
  PORT(
    twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_12_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_12_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_12_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_12_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_12_obj_twiddle_rsc_triosy_0_12_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_12_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_12_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_12_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_12_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_12_obj_twiddle_rsc_triosy_0_12_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_12_obj_twiddle_rsc_triosy_0_12_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_12_obj_iswt0 => twiddle_rsc_triosy_0_12_obj_iswt0,
      twiddle_rsc_triosy_0_12_obj_ld_core_sct => twiddle_rsc_triosy_0_12_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_13_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_13_obj IS
  PORT(
    twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_13_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_13_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_13_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_13_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_13_obj_twiddle_rsc_triosy_0_13_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_13_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_13_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_13_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_13_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_13_obj_twiddle_rsc_triosy_0_13_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_13_obj_twiddle_rsc_triosy_0_13_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_13_obj_iswt0 => twiddle_rsc_triosy_0_13_obj_iswt0,
      twiddle_rsc_triosy_0_13_obj_ld_core_sct => twiddle_rsc_triosy_0_13_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_14_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_14_obj IS
  PORT(
    twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_14_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_14_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_14_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_14_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_14_obj_twiddle_rsc_triosy_0_14_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_14_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_14_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_14_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_14_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_14_obj_twiddle_rsc_triosy_0_14_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_14_obj_twiddle_rsc_triosy_0_14_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_14_obj_iswt0 => twiddle_rsc_triosy_0_14_obj_iswt0,
      twiddle_rsc_triosy_0_14_obj_ld_core_sct => twiddle_rsc_triosy_0_14_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_triosy_0_15_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_triosy_0_15_obj IS
  PORT(
    twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    twiddle_rsc_triosy_0_15_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_twiddle_rsc_triosy_0_15_obj;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_triosy_0_15_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_triosy_0_15_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_15_obj_twiddle_rsc_triosy_0_15_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_15_obj_iswt0 : IN STD_LOGIC;
      twiddle_rsc_triosy_0_15_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  twiddle_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => twiddle_rsc_triosy_0_15_obj_ld_core_sct,
      lz => twiddle_rsc_triosy_0_15_lz
    );
  peaseNTT_core_twiddle_rsc_triosy_0_15_obj_twiddle_rsc_triosy_0_15_wait_ctrl_inst
      : peaseNTT_core_twiddle_rsc_triosy_0_15_obj_twiddle_rsc_triosy_0_15_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      twiddle_rsc_triosy_0_15_obj_iswt0 => twiddle_rsc_triosy_0_15_obj_iswt0,
      twiddle_rsc_triosy_0_15_obj_ld_core_sct => twiddle_rsc_triosy_0_15_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_r_rsc_triosy_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_r_rsc_triosy_obj IS
  PORT(
    r_rsc_triosy_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    r_rsc_triosy_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_r_rsc_triosy_obj;

ARCHITECTURE v29 OF peaseNTT_core_r_rsc_triosy_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL r_rsc_triosy_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_r_rsc_triosy_obj_r_rsc_triosy_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      r_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
      r_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  r_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => r_rsc_triosy_obj_ld_core_sct,
      lz => r_rsc_triosy_lz
    );
  peaseNTT_core_r_rsc_triosy_obj_r_rsc_triosy_wait_ctrl_inst : peaseNTT_core_r_rsc_triosy_obj_r_rsc_triosy_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      r_rsc_triosy_obj_iswt0 => r_rsc_triosy_obj_iswt0,
      r_rsc_triosy_obj_ld_core_sct => r_rsc_triosy_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_p_rsc_triosy_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_p_rsc_triosy_obj IS
  PORT(
    p_rsc_triosy_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    p_rsc_triosy_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_p_rsc_triosy_obj;

ARCHITECTURE v29 OF peaseNTT_core_p_rsc_triosy_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL p_rsc_triosy_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_p_rsc_triosy_obj_p_rsc_triosy_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      p_rsc_triosy_obj_iswt0 : IN STD_LOGIC;
      p_rsc_triosy_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  p_rsc_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => p_rsc_triosy_obj_ld_core_sct,
      lz => p_rsc_triosy_lz
    );
  peaseNTT_core_p_rsc_triosy_obj_p_rsc_triosy_wait_ctrl_inst : peaseNTT_core_p_rsc_triosy_obj_p_rsc_triosy_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      p_rsc_triosy_obj_iswt0 => p_rsc_triosy_obj_iswt0,
      p_rsc_triosy_obj_ld_core_sct => p_rsc_triosy_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_0_obj IS
  PORT(
    xt_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_0_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_0_obj_xt_rsc_triosy_0_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_0_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_0_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_0_obj_xt_rsc_triosy_0_0_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_0_obj_xt_rsc_triosy_0_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_0_obj_iswt0 => xt_rsc_triosy_0_0_obj_iswt0,
      xt_rsc_triosy_0_0_obj_ld_core_sct => xt_rsc_triosy_0_0_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_1_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_1_obj IS
  PORT(
    xt_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_1_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_1_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_1_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_1_obj_xt_rsc_triosy_0_1_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_1_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_1_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_1_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_1_obj_xt_rsc_triosy_0_1_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_1_obj_xt_rsc_triosy_0_1_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_1_obj_iswt0 => xt_rsc_triosy_0_1_obj_iswt0,
      xt_rsc_triosy_0_1_obj_ld_core_sct => xt_rsc_triosy_0_1_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_2_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_2_obj IS
  PORT(
    xt_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_2_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_2_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_2_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_2_obj_xt_rsc_triosy_0_2_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_2_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_2_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_2_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_2_obj_xt_rsc_triosy_0_2_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_2_obj_xt_rsc_triosy_0_2_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_2_obj_iswt0 => xt_rsc_triosy_0_2_obj_iswt0,
      xt_rsc_triosy_0_2_obj_ld_core_sct => xt_rsc_triosy_0_2_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_3_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_3_obj IS
  PORT(
    xt_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_3_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_3_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_3_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_3_obj_xt_rsc_triosy_0_3_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_3_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_3_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_3_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_3_obj_xt_rsc_triosy_0_3_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_3_obj_xt_rsc_triosy_0_3_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_3_obj_iswt0 => xt_rsc_triosy_0_3_obj_iswt0,
      xt_rsc_triosy_0_3_obj_ld_core_sct => xt_rsc_triosy_0_3_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_4_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_4_obj IS
  PORT(
    xt_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_4_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_4_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_4_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_4_obj_xt_rsc_triosy_0_4_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_4_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_4_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_4_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_4_obj_xt_rsc_triosy_0_4_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_4_obj_xt_rsc_triosy_0_4_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_4_obj_iswt0 => xt_rsc_triosy_0_4_obj_iswt0,
      xt_rsc_triosy_0_4_obj_ld_core_sct => xt_rsc_triosy_0_4_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_5_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_5_obj IS
  PORT(
    xt_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_5_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_5_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_5_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_5_obj_xt_rsc_triosy_0_5_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_5_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_5_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_5_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_5_obj_xt_rsc_triosy_0_5_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_5_obj_xt_rsc_triosy_0_5_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_5_obj_iswt0 => xt_rsc_triosy_0_5_obj_iswt0,
      xt_rsc_triosy_0_5_obj_ld_core_sct => xt_rsc_triosy_0_5_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_6_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_6_obj IS
  PORT(
    xt_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_6_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_6_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_6_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_6_obj_xt_rsc_triosy_0_6_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_6_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_6_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_6_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_6_obj_xt_rsc_triosy_0_6_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_6_obj_xt_rsc_triosy_0_6_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_6_obj_iswt0 => xt_rsc_triosy_0_6_obj_iswt0,
      xt_rsc_triosy_0_6_obj_ld_core_sct => xt_rsc_triosy_0_6_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_7_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_7_obj IS
  PORT(
    xt_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_7_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_7_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_7_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_7_obj_xt_rsc_triosy_0_7_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_7_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_7_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_7_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_7_obj_xt_rsc_triosy_0_7_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_7_obj_xt_rsc_triosy_0_7_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_7_obj_iswt0 => xt_rsc_triosy_0_7_obj_iswt0,
      xt_rsc_triosy_0_7_obj_ld_core_sct => xt_rsc_triosy_0_7_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_8_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_8_obj IS
  PORT(
    xt_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_8_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_8_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_8_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_8_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_8_obj_xt_rsc_triosy_0_8_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_8_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_8_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_8_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_8_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_8_obj_xt_rsc_triosy_0_8_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_8_obj_xt_rsc_triosy_0_8_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_8_obj_iswt0 => xt_rsc_triosy_0_8_obj_iswt0,
      xt_rsc_triosy_0_8_obj_ld_core_sct => xt_rsc_triosy_0_8_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_9_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_9_obj IS
  PORT(
    xt_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_9_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_9_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_9_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_9_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_9_obj_xt_rsc_triosy_0_9_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_9_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_9_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_9_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_9_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_9_obj_xt_rsc_triosy_0_9_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_9_obj_xt_rsc_triosy_0_9_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_9_obj_iswt0 => xt_rsc_triosy_0_9_obj_iswt0,
      xt_rsc_triosy_0_9_obj_ld_core_sct => xt_rsc_triosy_0_9_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_10_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_10_obj IS
  PORT(
    xt_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_10_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_10_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_10_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_10_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_10_obj_xt_rsc_triosy_0_10_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_10_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_10_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_10_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_10_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_10_obj_xt_rsc_triosy_0_10_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_10_obj_xt_rsc_triosy_0_10_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_10_obj_iswt0 => xt_rsc_triosy_0_10_obj_iswt0,
      xt_rsc_triosy_0_10_obj_ld_core_sct => xt_rsc_triosy_0_10_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_11_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_11_obj IS
  PORT(
    xt_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_11_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_11_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_11_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_11_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_11_obj_xt_rsc_triosy_0_11_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_11_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_11_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_11_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_11_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_11_obj_xt_rsc_triosy_0_11_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_11_obj_xt_rsc_triosy_0_11_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_11_obj_iswt0 => xt_rsc_triosy_0_11_obj_iswt0,
      xt_rsc_triosy_0_11_obj_ld_core_sct => xt_rsc_triosy_0_11_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_12_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_12_obj IS
  PORT(
    xt_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_12_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_12_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_12_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_12_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_12_obj_xt_rsc_triosy_0_12_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_12_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_12_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_12_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_12_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_12_obj_xt_rsc_triosy_0_12_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_12_obj_xt_rsc_triosy_0_12_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_12_obj_iswt0 => xt_rsc_triosy_0_12_obj_iswt0,
      xt_rsc_triosy_0_12_obj_ld_core_sct => xt_rsc_triosy_0_12_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_13_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_13_obj IS
  PORT(
    xt_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_13_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_13_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_13_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_13_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_13_obj_xt_rsc_triosy_0_13_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_13_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_13_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_13_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_13_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_13_obj_xt_rsc_triosy_0_13_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_13_obj_xt_rsc_triosy_0_13_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_13_obj_iswt0 => xt_rsc_triosy_0_13_obj_iswt0,
      xt_rsc_triosy_0_13_obj_ld_core_sct => xt_rsc_triosy_0_13_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_14_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_14_obj IS
  PORT(
    xt_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_14_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_14_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_14_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_14_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_14_obj_xt_rsc_triosy_0_14_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_14_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_14_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_14_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_14_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_14_obj_xt_rsc_triosy_0_14_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_14_obj_xt_rsc_triosy_0_14_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_14_obj_iswt0 => xt_rsc_triosy_0_14_obj_iswt0,
      xt_rsc_triosy_0_14_obj_ld_core_sct => xt_rsc_triosy_0_14_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_15_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_15_obj IS
  PORT(
    xt_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_15_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_15_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_15_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_15_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_15_obj_xt_rsc_triosy_0_15_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_15_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_15_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_15_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_15_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_15_obj_xt_rsc_triosy_0_15_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_15_obj_xt_rsc_triosy_0_15_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_15_obj_iswt0 => xt_rsc_triosy_0_15_obj_iswt0,
      xt_rsc_triosy_0_15_obj_ld_core_sct => xt_rsc_triosy_0_15_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_16_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_16_obj IS
  PORT(
    xt_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_16_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_16_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_16_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_16_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_16_obj_xt_rsc_triosy_0_16_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_16_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_16_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_16_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_16_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_16_obj_xt_rsc_triosy_0_16_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_16_obj_xt_rsc_triosy_0_16_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_16_obj_iswt0 => xt_rsc_triosy_0_16_obj_iswt0,
      xt_rsc_triosy_0_16_obj_ld_core_sct => xt_rsc_triosy_0_16_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_17_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_17_obj IS
  PORT(
    xt_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_17_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_17_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_17_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_17_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_17_obj_xt_rsc_triosy_0_17_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_17_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_17_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_17_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_17_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_17_obj_xt_rsc_triosy_0_17_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_17_obj_xt_rsc_triosy_0_17_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_17_obj_iswt0 => xt_rsc_triosy_0_17_obj_iswt0,
      xt_rsc_triosy_0_17_obj_ld_core_sct => xt_rsc_triosy_0_17_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_18_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_18_obj IS
  PORT(
    xt_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_18_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_18_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_18_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_18_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_18_obj_xt_rsc_triosy_0_18_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_18_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_18_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_18_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_18_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_18_obj_xt_rsc_triosy_0_18_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_18_obj_xt_rsc_triosy_0_18_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_18_obj_iswt0 => xt_rsc_triosy_0_18_obj_iswt0,
      xt_rsc_triosy_0_18_obj_ld_core_sct => xt_rsc_triosy_0_18_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_19_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_19_obj IS
  PORT(
    xt_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_19_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_19_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_19_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_19_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_19_obj_xt_rsc_triosy_0_19_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_19_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_19_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_19_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_19_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_19_obj_xt_rsc_triosy_0_19_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_19_obj_xt_rsc_triosy_0_19_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_19_obj_iswt0 => xt_rsc_triosy_0_19_obj_iswt0,
      xt_rsc_triosy_0_19_obj_ld_core_sct => xt_rsc_triosy_0_19_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_20_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_20_obj IS
  PORT(
    xt_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_20_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_20_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_20_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_20_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_20_obj_xt_rsc_triosy_0_20_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_20_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_20_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_20_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_20_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_20_obj_xt_rsc_triosy_0_20_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_20_obj_xt_rsc_triosy_0_20_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_20_obj_iswt0 => xt_rsc_triosy_0_20_obj_iswt0,
      xt_rsc_triosy_0_20_obj_ld_core_sct => xt_rsc_triosy_0_20_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_21_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_21_obj IS
  PORT(
    xt_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_21_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_21_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_21_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_21_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_21_obj_xt_rsc_triosy_0_21_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_21_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_21_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_21_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_21_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_21_obj_xt_rsc_triosy_0_21_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_21_obj_xt_rsc_triosy_0_21_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_21_obj_iswt0 => xt_rsc_triosy_0_21_obj_iswt0,
      xt_rsc_triosy_0_21_obj_ld_core_sct => xt_rsc_triosy_0_21_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_22_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_22_obj IS
  PORT(
    xt_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_22_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_22_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_22_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_22_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_22_obj_xt_rsc_triosy_0_22_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_22_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_22_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_22_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_22_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_22_obj_xt_rsc_triosy_0_22_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_22_obj_xt_rsc_triosy_0_22_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_22_obj_iswt0 => xt_rsc_triosy_0_22_obj_iswt0,
      xt_rsc_triosy_0_22_obj_ld_core_sct => xt_rsc_triosy_0_22_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_23_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_23_obj IS
  PORT(
    xt_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_23_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_23_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_23_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_23_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_23_obj_xt_rsc_triosy_0_23_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_23_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_23_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_23_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_23_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_23_obj_xt_rsc_triosy_0_23_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_23_obj_xt_rsc_triosy_0_23_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_23_obj_iswt0 => xt_rsc_triosy_0_23_obj_iswt0,
      xt_rsc_triosy_0_23_obj_ld_core_sct => xt_rsc_triosy_0_23_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_24_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_24_obj IS
  PORT(
    xt_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_24_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_24_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_24_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_24_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_24_obj_xt_rsc_triosy_0_24_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_24_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_24_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_24_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_24_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_24_obj_xt_rsc_triosy_0_24_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_24_obj_xt_rsc_triosy_0_24_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_24_obj_iswt0 => xt_rsc_triosy_0_24_obj_iswt0,
      xt_rsc_triosy_0_24_obj_ld_core_sct => xt_rsc_triosy_0_24_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_25_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_25_obj IS
  PORT(
    xt_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_25_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_25_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_25_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_25_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_25_obj_xt_rsc_triosy_0_25_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_25_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_25_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_25_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_25_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_25_obj_xt_rsc_triosy_0_25_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_25_obj_xt_rsc_triosy_0_25_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_25_obj_iswt0 => xt_rsc_triosy_0_25_obj_iswt0,
      xt_rsc_triosy_0_25_obj_ld_core_sct => xt_rsc_triosy_0_25_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_26_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_26_obj IS
  PORT(
    xt_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_26_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_26_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_26_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_26_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_26_obj_xt_rsc_triosy_0_26_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_26_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_26_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_26_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_26_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_26_obj_xt_rsc_triosy_0_26_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_26_obj_xt_rsc_triosy_0_26_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_26_obj_iswt0 => xt_rsc_triosy_0_26_obj_iswt0,
      xt_rsc_triosy_0_26_obj_ld_core_sct => xt_rsc_triosy_0_26_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_27_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_27_obj IS
  PORT(
    xt_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_27_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_27_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_27_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_27_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_27_obj_xt_rsc_triosy_0_27_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_27_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_27_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_27_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_27_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_27_obj_xt_rsc_triosy_0_27_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_27_obj_xt_rsc_triosy_0_27_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_27_obj_iswt0 => xt_rsc_triosy_0_27_obj_iswt0,
      xt_rsc_triosy_0_27_obj_ld_core_sct => xt_rsc_triosy_0_27_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_28_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_28_obj IS
  PORT(
    xt_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_28_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_28_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_28_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_28_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_28_obj_xt_rsc_triosy_0_28_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_28_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_28_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_28_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_28_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_28_obj_xt_rsc_triosy_0_28_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_28_obj_xt_rsc_triosy_0_28_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_28_obj_iswt0 => xt_rsc_triosy_0_28_obj_iswt0,
      xt_rsc_triosy_0_28_obj_ld_core_sct => xt_rsc_triosy_0_28_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_29_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_29_obj IS
  PORT(
    xt_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_29_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_29_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_29_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_29_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_29_obj_xt_rsc_triosy_0_29_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_29_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_29_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_29_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_29_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_29_obj_xt_rsc_triosy_0_29_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_29_obj_xt_rsc_triosy_0_29_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_29_obj_iswt0 => xt_rsc_triosy_0_29_obj_iswt0,
      xt_rsc_triosy_0_29_obj_ld_core_sct => xt_rsc_triosy_0_29_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_30_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_30_obj IS
  PORT(
    xt_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_30_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_30_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_30_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_30_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_30_obj_xt_rsc_triosy_0_30_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_30_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_30_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_30_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_30_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_30_obj_xt_rsc_triosy_0_30_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_30_obj_xt_rsc_triosy_0_30_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_30_obj_iswt0 => xt_rsc_triosy_0_30_obj_iswt0,
      xt_rsc_triosy_0_30_obj_ld_core_sct => xt_rsc_triosy_0_30_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_0_31_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_0_31_obj IS
  PORT(
    xt_rsc_triosy_0_31_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_0_31_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_0_31_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_0_31_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_0_31_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_0_31_obj_xt_rsc_triosy_0_31_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_31_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_0_31_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_0_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_0_31_obj_ld_core_sct,
      lz => xt_rsc_triosy_0_31_lz
    );
  peaseNTT_core_xt_rsc_triosy_0_31_obj_xt_rsc_triosy_0_31_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_0_31_obj_xt_rsc_triosy_0_31_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_0_31_obj_iswt0 => xt_rsc_triosy_0_31_obj_iswt0,
      xt_rsc_triosy_0_31_obj_ld_core_sct => xt_rsc_triosy_0_31_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_0_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_0_obj IS
  PORT(
    xt_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_0_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_0_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_0_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_0_obj_xt_rsc_triosy_1_0_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_0_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_0_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_0_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_0_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_0_obj_xt_rsc_triosy_1_0_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_0_obj_xt_rsc_triosy_1_0_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_0_obj_iswt0 => xt_rsc_triosy_1_0_obj_iswt0,
      xt_rsc_triosy_1_0_obj_ld_core_sct => xt_rsc_triosy_1_0_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_1_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_1_obj IS
  PORT(
    xt_rsc_triosy_1_1_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_1_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_1_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_1_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_1_obj_xt_rsc_triosy_1_1_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_1_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_1_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_1_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_1_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_1_obj_xt_rsc_triosy_1_1_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_1_obj_xt_rsc_triosy_1_1_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_1_obj_iswt0 => xt_rsc_triosy_1_1_obj_iswt0,
      xt_rsc_triosy_1_1_obj_ld_core_sct => xt_rsc_triosy_1_1_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_2_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_2_obj IS
  PORT(
    xt_rsc_triosy_1_2_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_2_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_2_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_2_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_2_obj_xt_rsc_triosy_1_2_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_2_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_2_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_2_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_2_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_2_obj_xt_rsc_triosy_1_2_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_2_obj_xt_rsc_triosy_1_2_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_2_obj_iswt0 => xt_rsc_triosy_1_2_obj_iswt0,
      xt_rsc_triosy_1_2_obj_ld_core_sct => xt_rsc_triosy_1_2_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_3_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_3_obj IS
  PORT(
    xt_rsc_triosy_1_3_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_3_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_3_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_3_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_3_obj_xt_rsc_triosy_1_3_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_3_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_3_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_3_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_3_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_3_obj_xt_rsc_triosy_1_3_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_3_obj_xt_rsc_triosy_1_3_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_3_obj_iswt0 => xt_rsc_triosy_1_3_obj_iswt0,
      xt_rsc_triosy_1_3_obj_ld_core_sct => xt_rsc_triosy_1_3_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_4_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_4_obj IS
  PORT(
    xt_rsc_triosy_1_4_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_4_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_4_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_4_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_4_obj_xt_rsc_triosy_1_4_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_4_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_4_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_4_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_4_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_4_obj_xt_rsc_triosy_1_4_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_4_obj_xt_rsc_triosy_1_4_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_4_obj_iswt0 => xt_rsc_triosy_1_4_obj_iswt0,
      xt_rsc_triosy_1_4_obj_ld_core_sct => xt_rsc_triosy_1_4_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_5_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_5_obj IS
  PORT(
    xt_rsc_triosy_1_5_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_5_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_5_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_5_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_5_obj_xt_rsc_triosy_1_5_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_5_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_5_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_5_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_5_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_5_obj_xt_rsc_triosy_1_5_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_5_obj_xt_rsc_triosy_1_5_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_5_obj_iswt0 => xt_rsc_triosy_1_5_obj_iswt0,
      xt_rsc_triosy_1_5_obj_ld_core_sct => xt_rsc_triosy_1_5_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_6_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_6_obj IS
  PORT(
    xt_rsc_triosy_1_6_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_6_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_6_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_6_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_6_obj_xt_rsc_triosy_1_6_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_6_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_6_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_6_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_6_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_6_obj_xt_rsc_triosy_1_6_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_6_obj_xt_rsc_triosy_1_6_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_6_obj_iswt0 => xt_rsc_triosy_1_6_obj_iswt0,
      xt_rsc_triosy_1_6_obj_ld_core_sct => xt_rsc_triosy_1_6_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_7_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_7_obj IS
  PORT(
    xt_rsc_triosy_1_7_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_7_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_7_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_7_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_7_obj_xt_rsc_triosy_1_7_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_7_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_7_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_7_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_7_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_7_obj_xt_rsc_triosy_1_7_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_7_obj_xt_rsc_triosy_1_7_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_7_obj_iswt0 => xt_rsc_triosy_1_7_obj_iswt0,
      xt_rsc_triosy_1_7_obj_ld_core_sct => xt_rsc_triosy_1_7_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_8_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_8_obj IS
  PORT(
    xt_rsc_triosy_1_8_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_8_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_8_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_8_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_8_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_8_obj_xt_rsc_triosy_1_8_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_8_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_8_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_8_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_8_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_8_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_8_obj_xt_rsc_triosy_1_8_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_8_obj_xt_rsc_triosy_1_8_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_8_obj_iswt0 => xt_rsc_triosy_1_8_obj_iswt0,
      xt_rsc_triosy_1_8_obj_ld_core_sct => xt_rsc_triosy_1_8_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_9_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_9_obj IS
  PORT(
    xt_rsc_triosy_1_9_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_9_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_9_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_9_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_9_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_9_obj_xt_rsc_triosy_1_9_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_9_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_9_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_9_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_9_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_9_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_9_obj_xt_rsc_triosy_1_9_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_9_obj_xt_rsc_triosy_1_9_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_9_obj_iswt0 => xt_rsc_triosy_1_9_obj_iswt0,
      xt_rsc_triosy_1_9_obj_ld_core_sct => xt_rsc_triosy_1_9_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_10_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_10_obj IS
  PORT(
    xt_rsc_triosy_1_10_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_10_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_10_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_10_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_10_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_10_obj_xt_rsc_triosy_1_10_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_10_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_10_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_10_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_10_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_10_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_10_obj_xt_rsc_triosy_1_10_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_10_obj_xt_rsc_triosy_1_10_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_10_obj_iswt0 => xt_rsc_triosy_1_10_obj_iswt0,
      xt_rsc_triosy_1_10_obj_ld_core_sct => xt_rsc_triosy_1_10_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_11_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_11_obj IS
  PORT(
    xt_rsc_triosy_1_11_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_11_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_11_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_11_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_11_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_11_obj_xt_rsc_triosy_1_11_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_11_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_11_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_11_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_11_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_11_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_11_obj_xt_rsc_triosy_1_11_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_11_obj_xt_rsc_triosy_1_11_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_11_obj_iswt0 => xt_rsc_triosy_1_11_obj_iswt0,
      xt_rsc_triosy_1_11_obj_ld_core_sct => xt_rsc_triosy_1_11_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_12_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_12_obj IS
  PORT(
    xt_rsc_triosy_1_12_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_12_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_12_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_12_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_12_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_12_obj_xt_rsc_triosy_1_12_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_12_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_12_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_12_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_12_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_12_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_12_obj_xt_rsc_triosy_1_12_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_12_obj_xt_rsc_triosy_1_12_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_12_obj_iswt0 => xt_rsc_triosy_1_12_obj_iswt0,
      xt_rsc_triosy_1_12_obj_ld_core_sct => xt_rsc_triosy_1_12_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_13_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_13_obj IS
  PORT(
    xt_rsc_triosy_1_13_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_13_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_13_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_13_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_13_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_13_obj_xt_rsc_triosy_1_13_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_13_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_13_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_13_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_13_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_13_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_13_obj_xt_rsc_triosy_1_13_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_13_obj_xt_rsc_triosy_1_13_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_13_obj_iswt0 => xt_rsc_triosy_1_13_obj_iswt0,
      xt_rsc_triosy_1_13_obj_ld_core_sct => xt_rsc_triosy_1_13_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_14_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_14_obj IS
  PORT(
    xt_rsc_triosy_1_14_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_14_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_14_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_14_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_14_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_14_obj_xt_rsc_triosy_1_14_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_14_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_14_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_14_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_14_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_14_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_14_obj_xt_rsc_triosy_1_14_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_14_obj_xt_rsc_triosy_1_14_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_14_obj_iswt0 => xt_rsc_triosy_1_14_obj_iswt0,
      xt_rsc_triosy_1_14_obj_ld_core_sct => xt_rsc_triosy_1_14_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_15_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_15_obj IS
  PORT(
    xt_rsc_triosy_1_15_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_15_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_15_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_15_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_15_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_15_obj_xt_rsc_triosy_1_15_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_15_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_15_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_15_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_15_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_15_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_15_obj_xt_rsc_triosy_1_15_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_15_obj_xt_rsc_triosy_1_15_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_15_obj_iswt0 => xt_rsc_triosy_1_15_obj_iswt0,
      xt_rsc_triosy_1_15_obj_ld_core_sct => xt_rsc_triosy_1_15_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_16_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_16_obj IS
  PORT(
    xt_rsc_triosy_1_16_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_16_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_16_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_16_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_16_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_16_obj_xt_rsc_triosy_1_16_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_16_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_16_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_16_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_16_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_16_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_16_obj_xt_rsc_triosy_1_16_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_16_obj_xt_rsc_triosy_1_16_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_16_obj_iswt0 => xt_rsc_triosy_1_16_obj_iswt0,
      xt_rsc_triosy_1_16_obj_ld_core_sct => xt_rsc_triosy_1_16_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_17_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_17_obj IS
  PORT(
    xt_rsc_triosy_1_17_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_17_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_17_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_17_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_17_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_17_obj_xt_rsc_triosy_1_17_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_17_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_17_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_17_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_17_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_17_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_17_obj_xt_rsc_triosy_1_17_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_17_obj_xt_rsc_triosy_1_17_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_17_obj_iswt0 => xt_rsc_triosy_1_17_obj_iswt0,
      xt_rsc_triosy_1_17_obj_ld_core_sct => xt_rsc_triosy_1_17_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_18_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_18_obj IS
  PORT(
    xt_rsc_triosy_1_18_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_18_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_18_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_18_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_18_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_18_obj_xt_rsc_triosy_1_18_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_18_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_18_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_18_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_18_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_18_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_18_obj_xt_rsc_triosy_1_18_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_18_obj_xt_rsc_triosy_1_18_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_18_obj_iswt0 => xt_rsc_triosy_1_18_obj_iswt0,
      xt_rsc_triosy_1_18_obj_ld_core_sct => xt_rsc_triosy_1_18_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_19_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_19_obj IS
  PORT(
    xt_rsc_triosy_1_19_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_19_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_19_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_19_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_19_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_19_obj_xt_rsc_triosy_1_19_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_19_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_19_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_19_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_19_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_19_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_19_obj_xt_rsc_triosy_1_19_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_19_obj_xt_rsc_triosy_1_19_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_19_obj_iswt0 => xt_rsc_triosy_1_19_obj_iswt0,
      xt_rsc_triosy_1_19_obj_ld_core_sct => xt_rsc_triosy_1_19_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_20_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_20_obj IS
  PORT(
    xt_rsc_triosy_1_20_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_20_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_20_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_20_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_20_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_20_obj_xt_rsc_triosy_1_20_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_20_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_20_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_20_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_20_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_20_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_20_obj_xt_rsc_triosy_1_20_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_20_obj_xt_rsc_triosy_1_20_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_20_obj_iswt0 => xt_rsc_triosy_1_20_obj_iswt0,
      xt_rsc_triosy_1_20_obj_ld_core_sct => xt_rsc_triosy_1_20_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_21_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_21_obj IS
  PORT(
    xt_rsc_triosy_1_21_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_21_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_21_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_21_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_21_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_21_obj_xt_rsc_triosy_1_21_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_21_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_21_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_21_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_21_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_21_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_21_obj_xt_rsc_triosy_1_21_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_21_obj_xt_rsc_triosy_1_21_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_21_obj_iswt0 => xt_rsc_triosy_1_21_obj_iswt0,
      xt_rsc_triosy_1_21_obj_ld_core_sct => xt_rsc_triosy_1_21_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_22_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_22_obj IS
  PORT(
    xt_rsc_triosy_1_22_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_22_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_22_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_22_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_22_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_22_obj_xt_rsc_triosy_1_22_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_22_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_22_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_22_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_22_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_22_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_22_obj_xt_rsc_triosy_1_22_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_22_obj_xt_rsc_triosy_1_22_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_22_obj_iswt0 => xt_rsc_triosy_1_22_obj_iswt0,
      xt_rsc_triosy_1_22_obj_ld_core_sct => xt_rsc_triosy_1_22_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_23_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_23_obj IS
  PORT(
    xt_rsc_triosy_1_23_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_23_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_23_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_23_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_23_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_23_obj_xt_rsc_triosy_1_23_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_23_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_23_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_23_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_23_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_23_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_23_obj_xt_rsc_triosy_1_23_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_23_obj_xt_rsc_triosy_1_23_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_23_obj_iswt0 => xt_rsc_triosy_1_23_obj_iswt0,
      xt_rsc_triosy_1_23_obj_ld_core_sct => xt_rsc_triosy_1_23_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_24_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_24_obj IS
  PORT(
    xt_rsc_triosy_1_24_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_24_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_24_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_24_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_24_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_24_obj_xt_rsc_triosy_1_24_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_24_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_24_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_24_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_24_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_24_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_24_obj_xt_rsc_triosy_1_24_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_24_obj_xt_rsc_triosy_1_24_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_24_obj_iswt0 => xt_rsc_triosy_1_24_obj_iswt0,
      xt_rsc_triosy_1_24_obj_ld_core_sct => xt_rsc_triosy_1_24_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_25_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_25_obj IS
  PORT(
    xt_rsc_triosy_1_25_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_25_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_25_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_25_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_25_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_25_obj_xt_rsc_triosy_1_25_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_25_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_25_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_25_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_25_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_25_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_25_obj_xt_rsc_triosy_1_25_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_25_obj_xt_rsc_triosy_1_25_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_25_obj_iswt0 => xt_rsc_triosy_1_25_obj_iswt0,
      xt_rsc_triosy_1_25_obj_ld_core_sct => xt_rsc_triosy_1_25_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_26_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_26_obj IS
  PORT(
    xt_rsc_triosy_1_26_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_26_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_26_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_26_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_26_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_26_obj_xt_rsc_triosy_1_26_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_26_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_26_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_26_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_26_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_26_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_26_obj_xt_rsc_triosy_1_26_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_26_obj_xt_rsc_triosy_1_26_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_26_obj_iswt0 => xt_rsc_triosy_1_26_obj_iswt0,
      xt_rsc_triosy_1_26_obj_ld_core_sct => xt_rsc_triosy_1_26_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_27_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_27_obj IS
  PORT(
    xt_rsc_triosy_1_27_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_27_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_27_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_27_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_27_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_27_obj_xt_rsc_triosy_1_27_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_27_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_27_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_27_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_27_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_27_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_27_obj_xt_rsc_triosy_1_27_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_27_obj_xt_rsc_triosy_1_27_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_27_obj_iswt0 => xt_rsc_triosy_1_27_obj_iswt0,
      xt_rsc_triosy_1_27_obj_ld_core_sct => xt_rsc_triosy_1_27_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_28_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_28_obj IS
  PORT(
    xt_rsc_triosy_1_28_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_28_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_28_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_28_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_28_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_28_obj_xt_rsc_triosy_1_28_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_28_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_28_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_28_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_28_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_28_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_28_obj_xt_rsc_triosy_1_28_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_28_obj_xt_rsc_triosy_1_28_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_28_obj_iswt0 => xt_rsc_triosy_1_28_obj_iswt0,
      xt_rsc_triosy_1_28_obj_ld_core_sct => xt_rsc_triosy_1_28_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_29_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_29_obj IS
  PORT(
    xt_rsc_triosy_1_29_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_29_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_29_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_29_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_29_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_29_obj_xt_rsc_triosy_1_29_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_29_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_29_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_29_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_29_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_29_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_29_obj_xt_rsc_triosy_1_29_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_29_obj_xt_rsc_triosy_1_29_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_29_obj_iswt0 => xt_rsc_triosy_1_29_obj_iswt0,
      xt_rsc_triosy_1_29_obj_ld_core_sct => xt_rsc_triosy_1_29_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_30_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_30_obj IS
  PORT(
    xt_rsc_triosy_1_30_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_30_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_30_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_30_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_30_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_30_obj_xt_rsc_triosy_1_30_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_30_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_30_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_30_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_30_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_30_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_30_obj_xt_rsc_triosy_1_30_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_30_obj_xt_rsc_triosy_1_30_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_30_obj_iswt0 => xt_rsc_triosy_1_30_obj_iswt0,
      xt_rsc_triosy_1_30_obj_ld_core_sct => xt_rsc_triosy_1_30_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_triosy_1_31_obj
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_triosy_1_31_obj IS
  PORT(
    xt_rsc_triosy_1_31_lz : OUT STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_triosy_1_31_obj_iswt0 : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_triosy_1_31_obj;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_triosy_1_31_obj IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL xt_rsc_triosy_1_31_obj_ld_core_sct : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_31_obj_xt_rsc_triosy_1_31_wait_ctrl
    PORT(
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_31_obj_iswt0 : IN STD_LOGIC;
      xt_rsc_triosy_1_31_obj_ld_core_sct : OUT STD_LOGIC
    );
  END COMPONENT;
BEGIN
  xt_rsc_triosy_1_31_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => xt_rsc_triosy_1_31_obj_ld_core_sct,
      lz => xt_rsc_triosy_1_31_lz
    );
  peaseNTT_core_xt_rsc_triosy_1_31_obj_xt_rsc_triosy_1_31_wait_ctrl_inst : peaseNTT_core_xt_rsc_triosy_1_31_obj_xt_rsc_triosy_1_31_wait_ctrl
    PORT MAP(
      core_wten => core_wten,
      xt_rsc_triosy_1_31_obj_iswt0 => xt_rsc_triosy_1_31_obj_iswt0,
      xt_rsc_triosy_1_31_obj_ld_core_sct => xt_rsc_triosy_1_31_obj_ld_core_sct
    );
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_15_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_15_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_15_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_15_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_15_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_15_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_15_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_15_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_15_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_15_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_15_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_15_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_15_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_15_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_15_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_15_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_15_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_15_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_15_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_15_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_15_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_15_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_15_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_15_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_15_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_15_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_15_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_15_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_15_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_15_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_15_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_15_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_15_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_15_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_15_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_15_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_15_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_15_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_15_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_15_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_15_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_15_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_15_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_15_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_15_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_15_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_15_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_15_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_15_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_15_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_15_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_15_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_15_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_15_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_15_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp_inst_twiddle_h_rsc_0_15_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp_inst_twiddle_h_rsc_0_15_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp_inst_twiddle_h_rsc_0_15_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp_inst_twiddle_h_rsc_0_15_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_15_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_15_i_AWID,
      AWADDR => twiddle_h_rsc_0_15_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_15_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_15_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_15_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_15_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_15_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_15_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_15_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_15_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_15_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_15_AWVALID,
      AWREADY => twiddle_h_rsc_0_15_AWREADY,
      WDATA => twiddle_h_rsc_0_15_i_WDATA,
      WSTRB => twiddle_h_rsc_0_15_i_WSTRB,
      WLAST => twiddle_h_rsc_0_15_WLAST,
      WUSER => twiddle_h_rsc_0_15_i_WUSER,
      WVALID => twiddle_h_rsc_0_15_WVALID,
      WREADY => twiddle_h_rsc_0_15_WREADY,
      BID => twiddle_h_rsc_0_15_i_BID,
      BRESP => twiddle_h_rsc_0_15_i_BRESP,
      BUSER => twiddle_h_rsc_0_15_i_BUSER,
      BVALID => twiddle_h_rsc_0_15_BVALID,
      BREADY => twiddle_h_rsc_0_15_BREADY,
      ARID => twiddle_h_rsc_0_15_i_ARID,
      ARADDR => twiddle_h_rsc_0_15_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_15_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_15_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_15_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_15_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_15_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_15_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_15_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_15_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_15_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_15_ARVALID,
      ARREADY => twiddle_h_rsc_0_15_ARREADY,
      RID => twiddle_h_rsc_0_15_i_RID,
      RDATA => twiddle_h_rsc_0_15_i_RDATA,
      RRESP => twiddle_h_rsc_0_15_i_RRESP,
      RLAST => twiddle_h_rsc_0_15_RLAST,
      RUSER => twiddle_h_rsc_0_15_i_RUSER,
      RVALID => twiddle_h_rsc_0_15_RVALID,
      RREADY => twiddle_h_rsc_0_15_RREADY,
      s_re => twiddle_h_rsc_0_15_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_15_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_15_i_s_waddr,
      s_din => twiddle_h_rsc_0_15_i_s_din_1,
      s_dout => twiddle_h_rsc_0_15_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_15_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_15_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_15_is_idle,
      tr_write_done => twiddle_h_rsc_0_15_tr_write_done,
      s_tdone => twiddle_h_rsc_0_15_s_tdone
    );
  twiddle_h_rsc_0_15_i_AWID(0) <= twiddle_h_rsc_0_15_AWID;
  twiddle_h_rsc_0_15_i_AWADDR <= twiddle_h_rsc_0_15_AWADDR;
  twiddle_h_rsc_0_15_i_AWLEN <= twiddle_h_rsc_0_15_AWLEN;
  twiddle_h_rsc_0_15_i_AWSIZE <= twiddle_h_rsc_0_15_AWSIZE;
  twiddle_h_rsc_0_15_i_AWBURST <= twiddle_h_rsc_0_15_AWBURST;
  twiddle_h_rsc_0_15_i_AWCACHE <= twiddle_h_rsc_0_15_AWCACHE;
  twiddle_h_rsc_0_15_i_AWPROT <= twiddle_h_rsc_0_15_AWPROT;
  twiddle_h_rsc_0_15_i_AWQOS <= twiddle_h_rsc_0_15_AWQOS;
  twiddle_h_rsc_0_15_i_AWREGION <= twiddle_h_rsc_0_15_AWREGION;
  twiddle_h_rsc_0_15_i_AWUSER(0) <= twiddle_h_rsc_0_15_AWUSER;
  twiddle_h_rsc_0_15_i_WDATA <= twiddle_h_rsc_0_15_WDATA;
  twiddle_h_rsc_0_15_i_WSTRB <= twiddle_h_rsc_0_15_WSTRB;
  twiddle_h_rsc_0_15_i_WUSER(0) <= twiddle_h_rsc_0_15_WUSER;
  twiddle_h_rsc_0_15_BID <= twiddle_h_rsc_0_15_i_BID(0);
  twiddle_h_rsc_0_15_BRESP <= twiddle_h_rsc_0_15_i_BRESP;
  twiddle_h_rsc_0_15_BUSER <= twiddle_h_rsc_0_15_i_BUSER(0);
  twiddle_h_rsc_0_15_i_ARID(0) <= twiddle_h_rsc_0_15_ARID;
  twiddle_h_rsc_0_15_i_ARADDR <= twiddle_h_rsc_0_15_ARADDR;
  twiddle_h_rsc_0_15_i_ARLEN <= twiddle_h_rsc_0_15_ARLEN;
  twiddle_h_rsc_0_15_i_ARSIZE <= twiddle_h_rsc_0_15_ARSIZE;
  twiddle_h_rsc_0_15_i_ARBURST <= twiddle_h_rsc_0_15_ARBURST;
  twiddle_h_rsc_0_15_i_ARCACHE <= twiddle_h_rsc_0_15_ARCACHE;
  twiddle_h_rsc_0_15_i_ARPROT <= twiddle_h_rsc_0_15_ARPROT;
  twiddle_h_rsc_0_15_i_ARQOS <= twiddle_h_rsc_0_15_ARQOS;
  twiddle_h_rsc_0_15_i_ARREGION <= twiddle_h_rsc_0_15_ARREGION;
  twiddle_h_rsc_0_15_i_ARUSER(0) <= twiddle_h_rsc_0_15_ARUSER;
  twiddle_h_rsc_0_15_RID <= twiddle_h_rsc_0_15_i_RID(0);
  twiddle_h_rsc_0_15_RDATA <= twiddle_h_rsc_0_15_i_RDATA;
  twiddle_h_rsc_0_15_RRESP <= twiddle_h_rsc_0_15_i_RRESP;
  twiddle_h_rsc_0_15_RUSER <= twiddle_h_rsc_0_15_i_RUSER(0);
  twiddle_h_rsc_0_15_i_s_raddr_1 <= twiddle_h_rsc_0_15_i_s_raddr;
  twiddle_h_rsc_0_15_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_15_i_s_din <= twiddle_h_rsc_0_15_i_s_din_1;
  twiddle_h_rsc_0_15_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_15_i_oswt => twiddle_h_rsc_0_15_i_oswt,
      twiddle_h_rsc_0_15_i_biwt => twiddle_h_rsc_0_15_i_biwt,
      twiddle_h_rsc_0_15_i_bdwt => twiddle_h_rsc_0_15_i_bdwt,
      twiddle_h_rsc_0_15_i_bcwt => twiddle_h_rsc_0_15_i_bcwt,
      twiddle_h_rsc_0_15_i_s_re_core_sct => twiddle_h_rsc_0_15_i_s_re_core_sct,
      twiddle_h_rsc_0_15_i_s_rrdy => twiddle_h_rsc_0_15_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_15_i_oswt => twiddle_h_rsc_0_15_i_oswt,
      twiddle_h_rsc_0_15_i_wen_comp => twiddle_h_rsc_0_15_i_wen_comp,
      twiddle_h_rsc_0_15_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp_inst_twiddle_h_rsc_0_15_i_s_raddr_core,
      twiddle_h_rsc_0_15_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp_inst_twiddle_h_rsc_0_15_i_s_din_mxwt,
      twiddle_h_rsc_0_15_i_biwt => twiddle_h_rsc_0_15_i_biwt,
      twiddle_h_rsc_0_15_i_bdwt => twiddle_h_rsc_0_15_i_bdwt,
      twiddle_h_rsc_0_15_i_bcwt => twiddle_h_rsc_0_15_i_bcwt,
      twiddle_h_rsc_0_15_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp_inst_twiddle_h_rsc_0_15_i_s_raddr,
      twiddle_h_rsc_0_15_i_s_raddr_core_sct => twiddle_h_rsc_0_15_i_s_re_core_sct,
      twiddle_h_rsc_0_15_i_s_din => peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp_inst_twiddle_h_rsc_0_15_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp_inst_twiddle_h_rsc_0_15_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_15_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_15_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp_inst_twiddle_h_rsc_0_15_i_s_din_mxwt;
  twiddle_h_rsc_0_15_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp_inst_twiddle_h_rsc_0_15_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_15_i_twiddle_h_rsc_0_15_wait_dp_inst_twiddle_h_rsc_0_15_i_s_din
      <= twiddle_h_rsc_0_15_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_14_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_14_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_14_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_14_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_14_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_14_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_14_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_14_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_14_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_14_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_14_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_14_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_14_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_14_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_14_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_14_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_14_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_14_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_14_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_14_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_14_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_14_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_14_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_14_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_14_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_14_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_14_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_14_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_14_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_14_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_14_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_14_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_14_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_14_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_14_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_14_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_14_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_14_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_14_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_14_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_14_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_14_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_14_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_14_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_14_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_14_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_14_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_14_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_14_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_14_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_14_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_14_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_14_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_14_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_14_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp_inst_twiddle_h_rsc_0_14_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp_inst_twiddle_h_rsc_0_14_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp_inst_twiddle_h_rsc_0_14_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp_inst_twiddle_h_rsc_0_14_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_14_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_14_i_AWID,
      AWADDR => twiddle_h_rsc_0_14_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_14_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_14_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_14_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_14_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_14_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_14_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_14_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_14_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_14_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_14_AWVALID,
      AWREADY => twiddle_h_rsc_0_14_AWREADY,
      WDATA => twiddle_h_rsc_0_14_i_WDATA,
      WSTRB => twiddle_h_rsc_0_14_i_WSTRB,
      WLAST => twiddle_h_rsc_0_14_WLAST,
      WUSER => twiddle_h_rsc_0_14_i_WUSER,
      WVALID => twiddle_h_rsc_0_14_WVALID,
      WREADY => twiddle_h_rsc_0_14_WREADY,
      BID => twiddle_h_rsc_0_14_i_BID,
      BRESP => twiddle_h_rsc_0_14_i_BRESP,
      BUSER => twiddle_h_rsc_0_14_i_BUSER,
      BVALID => twiddle_h_rsc_0_14_BVALID,
      BREADY => twiddle_h_rsc_0_14_BREADY,
      ARID => twiddle_h_rsc_0_14_i_ARID,
      ARADDR => twiddle_h_rsc_0_14_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_14_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_14_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_14_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_14_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_14_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_14_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_14_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_14_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_14_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_14_ARVALID,
      ARREADY => twiddle_h_rsc_0_14_ARREADY,
      RID => twiddle_h_rsc_0_14_i_RID,
      RDATA => twiddle_h_rsc_0_14_i_RDATA,
      RRESP => twiddle_h_rsc_0_14_i_RRESP,
      RLAST => twiddle_h_rsc_0_14_RLAST,
      RUSER => twiddle_h_rsc_0_14_i_RUSER,
      RVALID => twiddle_h_rsc_0_14_RVALID,
      RREADY => twiddle_h_rsc_0_14_RREADY,
      s_re => twiddle_h_rsc_0_14_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_14_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_14_i_s_waddr,
      s_din => twiddle_h_rsc_0_14_i_s_din_1,
      s_dout => twiddle_h_rsc_0_14_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_14_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_14_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_14_is_idle,
      tr_write_done => twiddle_h_rsc_0_14_tr_write_done,
      s_tdone => twiddle_h_rsc_0_14_s_tdone
    );
  twiddle_h_rsc_0_14_i_AWID(0) <= twiddle_h_rsc_0_14_AWID;
  twiddle_h_rsc_0_14_i_AWADDR <= twiddle_h_rsc_0_14_AWADDR;
  twiddle_h_rsc_0_14_i_AWLEN <= twiddle_h_rsc_0_14_AWLEN;
  twiddle_h_rsc_0_14_i_AWSIZE <= twiddle_h_rsc_0_14_AWSIZE;
  twiddle_h_rsc_0_14_i_AWBURST <= twiddle_h_rsc_0_14_AWBURST;
  twiddle_h_rsc_0_14_i_AWCACHE <= twiddle_h_rsc_0_14_AWCACHE;
  twiddle_h_rsc_0_14_i_AWPROT <= twiddle_h_rsc_0_14_AWPROT;
  twiddle_h_rsc_0_14_i_AWQOS <= twiddle_h_rsc_0_14_AWQOS;
  twiddle_h_rsc_0_14_i_AWREGION <= twiddle_h_rsc_0_14_AWREGION;
  twiddle_h_rsc_0_14_i_AWUSER(0) <= twiddle_h_rsc_0_14_AWUSER;
  twiddle_h_rsc_0_14_i_WDATA <= twiddle_h_rsc_0_14_WDATA;
  twiddle_h_rsc_0_14_i_WSTRB <= twiddle_h_rsc_0_14_WSTRB;
  twiddle_h_rsc_0_14_i_WUSER(0) <= twiddle_h_rsc_0_14_WUSER;
  twiddle_h_rsc_0_14_BID <= twiddle_h_rsc_0_14_i_BID(0);
  twiddle_h_rsc_0_14_BRESP <= twiddle_h_rsc_0_14_i_BRESP;
  twiddle_h_rsc_0_14_BUSER <= twiddle_h_rsc_0_14_i_BUSER(0);
  twiddle_h_rsc_0_14_i_ARID(0) <= twiddle_h_rsc_0_14_ARID;
  twiddle_h_rsc_0_14_i_ARADDR <= twiddle_h_rsc_0_14_ARADDR;
  twiddle_h_rsc_0_14_i_ARLEN <= twiddle_h_rsc_0_14_ARLEN;
  twiddle_h_rsc_0_14_i_ARSIZE <= twiddle_h_rsc_0_14_ARSIZE;
  twiddle_h_rsc_0_14_i_ARBURST <= twiddle_h_rsc_0_14_ARBURST;
  twiddle_h_rsc_0_14_i_ARCACHE <= twiddle_h_rsc_0_14_ARCACHE;
  twiddle_h_rsc_0_14_i_ARPROT <= twiddle_h_rsc_0_14_ARPROT;
  twiddle_h_rsc_0_14_i_ARQOS <= twiddle_h_rsc_0_14_ARQOS;
  twiddle_h_rsc_0_14_i_ARREGION <= twiddle_h_rsc_0_14_ARREGION;
  twiddle_h_rsc_0_14_i_ARUSER(0) <= twiddle_h_rsc_0_14_ARUSER;
  twiddle_h_rsc_0_14_RID <= twiddle_h_rsc_0_14_i_RID(0);
  twiddle_h_rsc_0_14_RDATA <= twiddle_h_rsc_0_14_i_RDATA;
  twiddle_h_rsc_0_14_RRESP <= twiddle_h_rsc_0_14_i_RRESP;
  twiddle_h_rsc_0_14_RUSER <= twiddle_h_rsc_0_14_i_RUSER(0);
  twiddle_h_rsc_0_14_i_s_raddr_1 <= twiddle_h_rsc_0_14_i_s_raddr;
  twiddle_h_rsc_0_14_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_14_i_s_din <= twiddle_h_rsc_0_14_i_s_din_1;
  twiddle_h_rsc_0_14_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_14_i_oswt => twiddle_h_rsc_0_14_i_oswt,
      twiddle_h_rsc_0_14_i_biwt => twiddle_h_rsc_0_14_i_biwt,
      twiddle_h_rsc_0_14_i_bdwt => twiddle_h_rsc_0_14_i_bdwt,
      twiddle_h_rsc_0_14_i_bcwt => twiddle_h_rsc_0_14_i_bcwt,
      twiddle_h_rsc_0_14_i_s_re_core_sct => twiddle_h_rsc_0_14_i_s_re_core_sct,
      twiddle_h_rsc_0_14_i_s_rrdy => twiddle_h_rsc_0_14_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_14_i_oswt => twiddle_h_rsc_0_14_i_oswt,
      twiddle_h_rsc_0_14_i_wen_comp => twiddle_h_rsc_0_14_i_wen_comp,
      twiddle_h_rsc_0_14_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp_inst_twiddle_h_rsc_0_14_i_s_raddr_core,
      twiddle_h_rsc_0_14_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp_inst_twiddle_h_rsc_0_14_i_s_din_mxwt,
      twiddle_h_rsc_0_14_i_biwt => twiddle_h_rsc_0_14_i_biwt,
      twiddle_h_rsc_0_14_i_bdwt => twiddle_h_rsc_0_14_i_bdwt,
      twiddle_h_rsc_0_14_i_bcwt => twiddle_h_rsc_0_14_i_bcwt,
      twiddle_h_rsc_0_14_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp_inst_twiddle_h_rsc_0_14_i_s_raddr,
      twiddle_h_rsc_0_14_i_s_raddr_core_sct => twiddle_h_rsc_0_14_i_s_re_core_sct,
      twiddle_h_rsc_0_14_i_s_din => peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp_inst_twiddle_h_rsc_0_14_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp_inst_twiddle_h_rsc_0_14_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_14_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_14_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp_inst_twiddle_h_rsc_0_14_i_s_din_mxwt;
  twiddle_h_rsc_0_14_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp_inst_twiddle_h_rsc_0_14_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_14_i_twiddle_h_rsc_0_14_wait_dp_inst_twiddle_h_rsc_0_14_i_s_din
      <= twiddle_h_rsc_0_14_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_13_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_13_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_13_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_13_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_13_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_13_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_13_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_13_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_13_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_13_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_13_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_13_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_13_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_13_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_13_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_13_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_13_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_13_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_13_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_13_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_13_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_13_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_13_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_13_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_13_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_13_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_13_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_13_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_13_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_13_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_13_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_13_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_13_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_13_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_13_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_13_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_13_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_13_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_13_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_13_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_13_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_13_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_13_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_13_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_13_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_13_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_13_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_13_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_13_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_13_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_13_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_13_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_13_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_13_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_13_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp_inst_twiddle_h_rsc_0_13_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp_inst_twiddle_h_rsc_0_13_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp_inst_twiddle_h_rsc_0_13_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp_inst_twiddle_h_rsc_0_13_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_13_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_13_i_AWID,
      AWADDR => twiddle_h_rsc_0_13_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_13_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_13_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_13_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_13_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_13_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_13_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_13_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_13_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_13_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_13_AWVALID,
      AWREADY => twiddle_h_rsc_0_13_AWREADY,
      WDATA => twiddle_h_rsc_0_13_i_WDATA,
      WSTRB => twiddle_h_rsc_0_13_i_WSTRB,
      WLAST => twiddle_h_rsc_0_13_WLAST,
      WUSER => twiddle_h_rsc_0_13_i_WUSER,
      WVALID => twiddle_h_rsc_0_13_WVALID,
      WREADY => twiddle_h_rsc_0_13_WREADY,
      BID => twiddle_h_rsc_0_13_i_BID,
      BRESP => twiddle_h_rsc_0_13_i_BRESP,
      BUSER => twiddle_h_rsc_0_13_i_BUSER,
      BVALID => twiddle_h_rsc_0_13_BVALID,
      BREADY => twiddle_h_rsc_0_13_BREADY,
      ARID => twiddle_h_rsc_0_13_i_ARID,
      ARADDR => twiddle_h_rsc_0_13_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_13_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_13_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_13_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_13_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_13_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_13_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_13_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_13_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_13_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_13_ARVALID,
      ARREADY => twiddle_h_rsc_0_13_ARREADY,
      RID => twiddle_h_rsc_0_13_i_RID,
      RDATA => twiddle_h_rsc_0_13_i_RDATA,
      RRESP => twiddle_h_rsc_0_13_i_RRESP,
      RLAST => twiddle_h_rsc_0_13_RLAST,
      RUSER => twiddle_h_rsc_0_13_i_RUSER,
      RVALID => twiddle_h_rsc_0_13_RVALID,
      RREADY => twiddle_h_rsc_0_13_RREADY,
      s_re => twiddle_h_rsc_0_13_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_13_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_13_i_s_waddr,
      s_din => twiddle_h_rsc_0_13_i_s_din_1,
      s_dout => twiddle_h_rsc_0_13_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_13_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_13_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_13_is_idle,
      tr_write_done => twiddle_h_rsc_0_13_tr_write_done,
      s_tdone => twiddle_h_rsc_0_13_s_tdone
    );
  twiddle_h_rsc_0_13_i_AWID(0) <= twiddle_h_rsc_0_13_AWID;
  twiddle_h_rsc_0_13_i_AWADDR <= twiddle_h_rsc_0_13_AWADDR;
  twiddle_h_rsc_0_13_i_AWLEN <= twiddle_h_rsc_0_13_AWLEN;
  twiddle_h_rsc_0_13_i_AWSIZE <= twiddle_h_rsc_0_13_AWSIZE;
  twiddle_h_rsc_0_13_i_AWBURST <= twiddle_h_rsc_0_13_AWBURST;
  twiddle_h_rsc_0_13_i_AWCACHE <= twiddle_h_rsc_0_13_AWCACHE;
  twiddle_h_rsc_0_13_i_AWPROT <= twiddle_h_rsc_0_13_AWPROT;
  twiddle_h_rsc_0_13_i_AWQOS <= twiddle_h_rsc_0_13_AWQOS;
  twiddle_h_rsc_0_13_i_AWREGION <= twiddle_h_rsc_0_13_AWREGION;
  twiddle_h_rsc_0_13_i_AWUSER(0) <= twiddle_h_rsc_0_13_AWUSER;
  twiddle_h_rsc_0_13_i_WDATA <= twiddle_h_rsc_0_13_WDATA;
  twiddle_h_rsc_0_13_i_WSTRB <= twiddle_h_rsc_0_13_WSTRB;
  twiddle_h_rsc_0_13_i_WUSER(0) <= twiddle_h_rsc_0_13_WUSER;
  twiddle_h_rsc_0_13_BID <= twiddle_h_rsc_0_13_i_BID(0);
  twiddle_h_rsc_0_13_BRESP <= twiddle_h_rsc_0_13_i_BRESP;
  twiddle_h_rsc_0_13_BUSER <= twiddle_h_rsc_0_13_i_BUSER(0);
  twiddle_h_rsc_0_13_i_ARID(0) <= twiddle_h_rsc_0_13_ARID;
  twiddle_h_rsc_0_13_i_ARADDR <= twiddle_h_rsc_0_13_ARADDR;
  twiddle_h_rsc_0_13_i_ARLEN <= twiddle_h_rsc_0_13_ARLEN;
  twiddle_h_rsc_0_13_i_ARSIZE <= twiddle_h_rsc_0_13_ARSIZE;
  twiddle_h_rsc_0_13_i_ARBURST <= twiddle_h_rsc_0_13_ARBURST;
  twiddle_h_rsc_0_13_i_ARCACHE <= twiddle_h_rsc_0_13_ARCACHE;
  twiddle_h_rsc_0_13_i_ARPROT <= twiddle_h_rsc_0_13_ARPROT;
  twiddle_h_rsc_0_13_i_ARQOS <= twiddle_h_rsc_0_13_ARQOS;
  twiddle_h_rsc_0_13_i_ARREGION <= twiddle_h_rsc_0_13_ARREGION;
  twiddle_h_rsc_0_13_i_ARUSER(0) <= twiddle_h_rsc_0_13_ARUSER;
  twiddle_h_rsc_0_13_RID <= twiddle_h_rsc_0_13_i_RID(0);
  twiddle_h_rsc_0_13_RDATA <= twiddle_h_rsc_0_13_i_RDATA;
  twiddle_h_rsc_0_13_RRESP <= twiddle_h_rsc_0_13_i_RRESP;
  twiddle_h_rsc_0_13_RUSER <= twiddle_h_rsc_0_13_i_RUSER(0);
  twiddle_h_rsc_0_13_i_s_raddr_1 <= twiddle_h_rsc_0_13_i_s_raddr;
  twiddle_h_rsc_0_13_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_13_i_s_din <= twiddle_h_rsc_0_13_i_s_din_1;
  twiddle_h_rsc_0_13_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_13_i_oswt => twiddle_h_rsc_0_13_i_oswt,
      twiddle_h_rsc_0_13_i_biwt => twiddle_h_rsc_0_13_i_biwt,
      twiddle_h_rsc_0_13_i_bdwt => twiddle_h_rsc_0_13_i_bdwt,
      twiddle_h_rsc_0_13_i_bcwt => twiddle_h_rsc_0_13_i_bcwt,
      twiddle_h_rsc_0_13_i_s_re_core_sct => twiddle_h_rsc_0_13_i_s_re_core_sct,
      twiddle_h_rsc_0_13_i_s_rrdy => twiddle_h_rsc_0_13_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_13_i_oswt => twiddle_h_rsc_0_13_i_oswt,
      twiddle_h_rsc_0_13_i_wen_comp => twiddle_h_rsc_0_13_i_wen_comp,
      twiddle_h_rsc_0_13_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp_inst_twiddle_h_rsc_0_13_i_s_raddr_core,
      twiddle_h_rsc_0_13_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp_inst_twiddle_h_rsc_0_13_i_s_din_mxwt,
      twiddle_h_rsc_0_13_i_biwt => twiddle_h_rsc_0_13_i_biwt,
      twiddle_h_rsc_0_13_i_bdwt => twiddle_h_rsc_0_13_i_bdwt,
      twiddle_h_rsc_0_13_i_bcwt => twiddle_h_rsc_0_13_i_bcwt,
      twiddle_h_rsc_0_13_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp_inst_twiddle_h_rsc_0_13_i_s_raddr,
      twiddle_h_rsc_0_13_i_s_raddr_core_sct => twiddle_h_rsc_0_13_i_s_re_core_sct,
      twiddle_h_rsc_0_13_i_s_din => peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp_inst_twiddle_h_rsc_0_13_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp_inst_twiddle_h_rsc_0_13_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_13_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_13_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp_inst_twiddle_h_rsc_0_13_i_s_din_mxwt;
  twiddle_h_rsc_0_13_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp_inst_twiddle_h_rsc_0_13_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_13_i_twiddle_h_rsc_0_13_wait_dp_inst_twiddle_h_rsc_0_13_i_s_din
      <= twiddle_h_rsc_0_13_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_12_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_12_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_12_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_12_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_12_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_12_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_12_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_12_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_12_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_12_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_12_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_12_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_12_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_12_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_12_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_12_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_12_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_12_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_12_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_12_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_12_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_12_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_12_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_12_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_12_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_12_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_12_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_12_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_12_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_12_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_12_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_12_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_12_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_12_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_12_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_12_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_12_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_12_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_12_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_12_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_12_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_12_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_12_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_12_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_12_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_12_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_12_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_12_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_12_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_12_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_12_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_12_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_12_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_12_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_12_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp_inst_twiddle_h_rsc_0_12_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp_inst_twiddle_h_rsc_0_12_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp_inst_twiddle_h_rsc_0_12_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp_inst_twiddle_h_rsc_0_12_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_12_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_12_i_AWID,
      AWADDR => twiddle_h_rsc_0_12_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_12_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_12_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_12_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_12_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_12_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_12_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_12_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_12_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_12_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_12_AWVALID,
      AWREADY => twiddle_h_rsc_0_12_AWREADY,
      WDATA => twiddle_h_rsc_0_12_i_WDATA,
      WSTRB => twiddle_h_rsc_0_12_i_WSTRB,
      WLAST => twiddle_h_rsc_0_12_WLAST,
      WUSER => twiddle_h_rsc_0_12_i_WUSER,
      WVALID => twiddle_h_rsc_0_12_WVALID,
      WREADY => twiddle_h_rsc_0_12_WREADY,
      BID => twiddle_h_rsc_0_12_i_BID,
      BRESP => twiddle_h_rsc_0_12_i_BRESP,
      BUSER => twiddle_h_rsc_0_12_i_BUSER,
      BVALID => twiddle_h_rsc_0_12_BVALID,
      BREADY => twiddle_h_rsc_0_12_BREADY,
      ARID => twiddle_h_rsc_0_12_i_ARID,
      ARADDR => twiddle_h_rsc_0_12_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_12_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_12_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_12_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_12_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_12_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_12_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_12_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_12_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_12_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_12_ARVALID,
      ARREADY => twiddle_h_rsc_0_12_ARREADY,
      RID => twiddle_h_rsc_0_12_i_RID,
      RDATA => twiddle_h_rsc_0_12_i_RDATA,
      RRESP => twiddle_h_rsc_0_12_i_RRESP,
      RLAST => twiddle_h_rsc_0_12_RLAST,
      RUSER => twiddle_h_rsc_0_12_i_RUSER,
      RVALID => twiddle_h_rsc_0_12_RVALID,
      RREADY => twiddle_h_rsc_0_12_RREADY,
      s_re => twiddle_h_rsc_0_12_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_12_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_12_i_s_waddr,
      s_din => twiddle_h_rsc_0_12_i_s_din_1,
      s_dout => twiddle_h_rsc_0_12_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_12_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_12_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_12_is_idle,
      tr_write_done => twiddle_h_rsc_0_12_tr_write_done,
      s_tdone => twiddle_h_rsc_0_12_s_tdone
    );
  twiddle_h_rsc_0_12_i_AWID(0) <= twiddle_h_rsc_0_12_AWID;
  twiddle_h_rsc_0_12_i_AWADDR <= twiddle_h_rsc_0_12_AWADDR;
  twiddle_h_rsc_0_12_i_AWLEN <= twiddle_h_rsc_0_12_AWLEN;
  twiddle_h_rsc_0_12_i_AWSIZE <= twiddle_h_rsc_0_12_AWSIZE;
  twiddle_h_rsc_0_12_i_AWBURST <= twiddle_h_rsc_0_12_AWBURST;
  twiddle_h_rsc_0_12_i_AWCACHE <= twiddle_h_rsc_0_12_AWCACHE;
  twiddle_h_rsc_0_12_i_AWPROT <= twiddle_h_rsc_0_12_AWPROT;
  twiddle_h_rsc_0_12_i_AWQOS <= twiddle_h_rsc_0_12_AWQOS;
  twiddle_h_rsc_0_12_i_AWREGION <= twiddle_h_rsc_0_12_AWREGION;
  twiddle_h_rsc_0_12_i_AWUSER(0) <= twiddle_h_rsc_0_12_AWUSER;
  twiddle_h_rsc_0_12_i_WDATA <= twiddle_h_rsc_0_12_WDATA;
  twiddle_h_rsc_0_12_i_WSTRB <= twiddle_h_rsc_0_12_WSTRB;
  twiddle_h_rsc_0_12_i_WUSER(0) <= twiddle_h_rsc_0_12_WUSER;
  twiddle_h_rsc_0_12_BID <= twiddle_h_rsc_0_12_i_BID(0);
  twiddle_h_rsc_0_12_BRESP <= twiddle_h_rsc_0_12_i_BRESP;
  twiddle_h_rsc_0_12_BUSER <= twiddle_h_rsc_0_12_i_BUSER(0);
  twiddle_h_rsc_0_12_i_ARID(0) <= twiddle_h_rsc_0_12_ARID;
  twiddle_h_rsc_0_12_i_ARADDR <= twiddle_h_rsc_0_12_ARADDR;
  twiddle_h_rsc_0_12_i_ARLEN <= twiddle_h_rsc_0_12_ARLEN;
  twiddle_h_rsc_0_12_i_ARSIZE <= twiddle_h_rsc_0_12_ARSIZE;
  twiddle_h_rsc_0_12_i_ARBURST <= twiddle_h_rsc_0_12_ARBURST;
  twiddle_h_rsc_0_12_i_ARCACHE <= twiddle_h_rsc_0_12_ARCACHE;
  twiddle_h_rsc_0_12_i_ARPROT <= twiddle_h_rsc_0_12_ARPROT;
  twiddle_h_rsc_0_12_i_ARQOS <= twiddle_h_rsc_0_12_ARQOS;
  twiddle_h_rsc_0_12_i_ARREGION <= twiddle_h_rsc_0_12_ARREGION;
  twiddle_h_rsc_0_12_i_ARUSER(0) <= twiddle_h_rsc_0_12_ARUSER;
  twiddle_h_rsc_0_12_RID <= twiddle_h_rsc_0_12_i_RID(0);
  twiddle_h_rsc_0_12_RDATA <= twiddle_h_rsc_0_12_i_RDATA;
  twiddle_h_rsc_0_12_RRESP <= twiddle_h_rsc_0_12_i_RRESP;
  twiddle_h_rsc_0_12_RUSER <= twiddle_h_rsc_0_12_i_RUSER(0);
  twiddle_h_rsc_0_12_i_s_raddr_1 <= twiddle_h_rsc_0_12_i_s_raddr;
  twiddle_h_rsc_0_12_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_12_i_s_din <= twiddle_h_rsc_0_12_i_s_din_1;
  twiddle_h_rsc_0_12_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_12_i_oswt => twiddle_h_rsc_0_12_i_oswt,
      twiddle_h_rsc_0_12_i_biwt => twiddle_h_rsc_0_12_i_biwt,
      twiddle_h_rsc_0_12_i_bdwt => twiddle_h_rsc_0_12_i_bdwt,
      twiddle_h_rsc_0_12_i_bcwt => twiddle_h_rsc_0_12_i_bcwt,
      twiddle_h_rsc_0_12_i_s_re_core_sct => twiddle_h_rsc_0_12_i_s_re_core_sct,
      twiddle_h_rsc_0_12_i_s_rrdy => twiddle_h_rsc_0_12_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_12_i_oswt => twiddle_h_rsc_0_12_i_oswt,
      twiddle_h_rsc_0_12_i_wen_comp => twiddle_h_rsc_0_12_i_wen_comp,
      twiddle_h_rsc_0_12_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp_inst_twiddle_h_rsc_0_12_i_s_raddr_core,
      twiddle_h_rsc_0_12_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp_inst_twiddle_h_rsc_0_12_i_s_din_mxwt,
      twiddle_h_rsc_0_12_i_biwt => twiddle_h_rsc_0_12_i_biwt,
      twiddle_h_rsc_0_12_i_bdwt => twiddle_h_rsc_0_12_i_bdwt,
      twiddle_h_rsc_0_12_i_bcwt => twiddle_h_rsc_0_12_i_bcwt,
      twiddle_h_rsc_0_12_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp_inst_twiddle_h_rsc_0_12_i_s_raddr,
      twiddle_h_rsc_0_12_i_s_raddr_core_sct => twiddle_h_rsc_0_12_i_s_re_core_sct,
      twiddle_h_rsc_0_12_i_s_din => peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp_inst_twiddle_h_rsc_0_12_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp_inst_twiddle_h_rsc_0_12_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_12_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_12_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp_inst_twiddle_h_rsc_0_12_i_s_din_mxwt;
  twiddle_h_rsc_0_12_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp_inst_twiddle_h_rsc_0_12_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_12_i_twiddle_h_rsc_0_12_wait_dp_inst_twiddle_h_rsc_0_12_i_s_din
      <= twiddle_h_rsc_0_12_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_11_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_11_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_11_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_11_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_11_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_11_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_11_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_11_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_11_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_11_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_11_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_11_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_11_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_11_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_11_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_11_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_11_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_11_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_11_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_11_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_11_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_11_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_11_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_11_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_11_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_11_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_11_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_11_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_11_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_11_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_11_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_11_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_11_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_11_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_11_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_11_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_11_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_11_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_11_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_11_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_11_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_11_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_11_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_11_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_11_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_11_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_11_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_11_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_11_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_11_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_11_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_11_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_11_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_11_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_11_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp_inst_twiddle_h_rsc_0_11_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp_inst_twiddle_h_rsc_0_11_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp_inst_twiddle_h_rsc_0_11_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp_inst_twiddle_h_rsc_0_11_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_11_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_11_i_AWID,
      AWADDR => twiddle_h_rsc_0_11_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_11_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_11_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_11_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_11_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_11_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_11_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_11_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_11_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_11_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_11_AWVALID,
      AWREADY => twiddle_h_rsc_0_11_AWREADY,
      WDATA => twiddle_h_rsc_0_11_i_WDATA,
      WSTRB => twiddle_h_rsc_0_11_i_WSTRB,
      WLAST => twiddle_h_rsc_0_11_WLAST,
      WUSER => twiddle_h_rsc_0_11_i_WUSER,
      WVALID => twiddle_h_rsc_0_11_WVALID,
      WREADY => twiddle_h_rsc_0_11_WREADY,
      BID => twiddle_h_rsc_0_11_i_BID,
      BRESP => twiddle_h_rsc_0_11_i_BRESP,
      BUSER => twiddle_h_rsc_0_11_i_BUSER,
      BVALID => twiddle_h_rsc_0_11_BVALID,
      BREADY => twiddle_h_rsc_0_11_BREADY,
      ARID => twiddle_h_rsc_0_11_i_ARID,
      ARADDR => twiddle_h_rsc_0_11_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_11_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_11_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_11_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_11_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_11_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_11_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_11_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_11_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_11_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_11_ARVALID,
      ARREADY => twiddle_h_rsc_0_11_ARREADY,
      RID => twiddle_h_rsc_0_11_i_RID,
      RDATA => twiddle_h_rsc_0_11_i_RDATA,
      RRESP => twiddle_h_rsc_0_11_i_RRESP,
      RLAST => twiddle_h_rsc_0_11_RLAST,
      RUSER => twiddle_h_rsc_0_11_i_RUSER,
      RVALID => twiddle_h_rsc_0_11_RVALID,
      RREADY => twiddle_h_rsc_0_11_RREADY,
      s_re => twiddle_h_rsc_0_11_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_11_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_11_i_s_waddr,
      s_din => twiddle_h_rsc_0_11_i_s_din_1,
      s_dout => twiddle_h_rsc_0_11_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_11_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_11_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_11_is_idle,
      tr_write_done => twiddle_h_rsc_0_11_tr_write_done,
      s_tdone => twiddle_h_rsc_0_11_s_tdone
    );
  twiddle_h_rsc_0_11_i_AWID(0) <= twiddle_h_rsc_0_11_AWID;
  twiddle_h_rsc_0_11_i_AWADDR <= twiddle_h_rsc_0_11_AWADDR;
  twiddle_h_rsc_0_11_i_AWLEN <= twiddle_h_rsc_0_11_AWLEN;
  twiddle_h_rsc_0_11_i_AWSIZE <= twiddle_h_rsc_0_11_AWSIZE;
  twiddle_h_rsc_0_11_i_AWBURST <= twiddle_h_rsc_0_11_AWBURST;
  twiddle_h_rsc_0_11_i_AWCACHE <= twiddle_h_rsc_0_11_AWCACHE;
  twiddle_h_rsc_0_11_i_AWPROT <= twiddle_h_rsc_0_11_AWPROT;
  twiddle_h_rsc_0_11_i_AWQOS <= twiddle_h_rsc_0_11_AWQOS;
  twiddle_h_rsc_0_11_i_AWREGION <= twiddle_h_rsc_0_11_AWREGION;
  twiddle_h_rsc_0_11_i_AWUSER(0) <= twiddle_h_rsc_0_11_AWUSER;
  twiddle_h_rsc_0_11_i_WDATA <= twiddle_h_rsc_0_11_WDATA;
  twiddle_h_rsc_0_11_i_WSTRB <= twiddle_h_rsc_0_11_WSTRB;
  twiddle_h_rsc_0_11_i_WUSER(0) <= twiddle_h_rsc_0_11_WUSER;
  twiddle_h_rsc_0_11_BID <= twiddle_h_rsc_0_11_i_BID(0);
  twiddle_h_rsc_0_11_BRESP <= twiddle_h_rsc_0_11_i_BRESP;
  twiddle_h_rsc_0_11_BUSER <= twiddle_h_rsc_0_11_i_BUSER(0);
  twiddle_h_rsc_0_11_i_ARID(0) <= twiddle_h_rsc_0_11_ARID;
  twiddle_h_rsc_0_11_i_ARADDR <= twiddle_h_rsc_0_11_ARADDR;
  twiddle_h_rsc_0_11_i_ARLEN <= twiddle_h_rsc_0_11_ARLEN;
  twiddle_h_rsc_0_11_i_ARSIZE <= twiddle_h_rsc_0_11_ARSIZE;
  twiddle_h_rsc_0_11_i_ARBURST <= twiddle_h_rsc_0_11_ARBURST;
  twiddle_h_rsc_0_11_i_ARCACHE <= twiddle_h_rsc_0_11_ARCACHE;
  twiddle_h_rsc_0_11_i_ARPROT <= twiddle_h_rsc_0_11_ARPROT;
  twiddle_h_rsc_0_11_i_ARQOS <= twiddle_h_rsc_0_11_ARQOS;
  twiddle_h_rsc_0_11_i_ARREGION <= twiddle_h_rsc_0_11_ARREGION;
  twiddle_h_rsc_0_11_i_ARUSER(0) <= twiddle_h_rsc_0_11_ARUSER;
  twiddle_h_rsc_0_11_RID <= twiddle_h_rsc_0_11_i_RID(0);
  twiddle_h_rsc_0_11_RDATA <= twiddle_h_rsc_0_11_i_RDATA;
  twiddle_h_rsc_0_11_RRESP <= twiddle_h_rsc_0_11_i_RRESP;
  twiddle_h_rsc_0_11_RUSER <= twiddle_h_rsc_0_11_i_RUSER(0);
  twiddle_h_rsc_0_11_i_s_raddr_1 <= twiddle_h_rsc_0_11_i_s_raddr;
  twiddle_h_rsc_0_11_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_11_i_s_din <= twiddle_h_rsc_0_11_i_s_din_1;
  twiddle_h_rsc_0_11_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_11_i_oswt => twiddle_h_rsc_0_11_i_oswt,
      twiddle_h_rsc_0_11_i_biwt => twiddle_h_rsc_0_11_i_biwt,
      twiddle_h_rsc_0_11_i_bdwt => twiddle_h_rsc_0_11_i_bdwt,
      twiddle_h_rsc_0_11_i_bcwt => twiddle_h_rsc_0_11_i_bcwt,
      twiddle_h_rsc_0_11_i_s_re_core_sct => twiddle_h_rsc_0_11_i_s_re_core_sct,
      twiddle_h_rsc_0_11_i_s_rrdy => twiddle_h_rsc_0_11_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_11_i_oswt => twiddle_h_rsc_0_11_i_oswt,
      twiddle_h_rsc_0_11_i_wen_comp => twiddle_h_rsc_0_11_i_wen_comp,
      twiddle_h_rsc_0_11_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp_inst_twiddle_h_rsc_0_11_i_s_raddr_core,
      twiddle_h_rsc_0_11_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp_inst_twiddle_h_rsc_0_11_i_s_din_mxwt,
      twiddle_h_rsc_0_11_i_biwt => twiddle_h_rsc_0_11_i_biwt,
      twiddle_h_rsc_0_11_i_bdwt => twiddle_h_rsc_0_11_i_bdwt,
      twiddle_h_rsc_0_11_i_bcwt => twiddle_h_rsc_0_11_i_bcwt,
      twiddle_h_rsc_0_11_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp_inst_twiddle_h_rsc_0_11_i_s_raddr,
      twiddle_h_rsc_0_11_i_s_raddr_core_sct => twiddle_h_rsc_0_11_i_s_re_core_sct,
      twiddle_h_rsc_0_11_i_s_din => peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp_inst_twiddle_h_rsc_0_11_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp_inst_twiddle_h_rsc_0_11_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_11_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_11_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp_inst_twiddle_h_rsc_0_11_i_s_din_mxwt;
  twiddle_h_rsc_0_11_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp_inst_twiddle_h_rsc_0_11_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_11_i_twiddle_h_rsc_0_11_wait_dp_inst_twiddle_h_rsc_0_11_i_s_din
      <= twiddle_h_rsc_0_11_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_10_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_10_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_10_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_10_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_10_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_10_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_10_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_10_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_10_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_10_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_10_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_10_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_10_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_10_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_10_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_10_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_10_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_10_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_10_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_10_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_10_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_10_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_10_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_10_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_10_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_10_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_10_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_10_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_10_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_10_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_10_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_10_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_10_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_10_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_10_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_10_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_10_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_10_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_10_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_10_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_10_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_10_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_10_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_10_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_10_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_10_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_10_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_10_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_10_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_10_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_10_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_10_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_10_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_10_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_10_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp_inst_twiddle_h_rsc_0_10_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp_inst_twiddle_h_rsc_0_10_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp_inst_twiddle_h_rsc_0_10_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp_inst_twiddle_h_rsc_0_10_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_10_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_10_i_AWID,
      AWADDR => twiddle_h_rsc_0_10_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_10_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_10_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_10_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_10_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_10_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_10_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_10_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_10_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_10_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_10_AWVALID,
      AWREADY => twiddle_h_rsc_0_10_AWREADY,
      WDATA => twiddle_h_rsc_0_10_i_WDATA,
      WSTRB => twiddle_h_rsc_0_10_i_WSTRB,
      WLAST => twiddle_h_rsc_0_10_WLAST,
      WUSER => twiddle_h_rsc_0_10_i_WUSER,
      WVALID => twiddle_h_rsc_0_10_WVALID,
      WREADY => twiddle_h_rsc_0_10_WREADY,
      BID => twiddle_h_rsc_0_10_i_BID,
      BRESP => twiddle_h_rsc_0_10_i_BRESP,
      BUSER => twiddle_h_rsc_0_10_i_BUSER,
      BVALID => twiddle_h_rsc_0_10_BVALID,
      BREADY => twiddle_h_rsc_0_10_BREADY,
      ARID => twiddle_h_rsc_0_10_i_ARID,
      ARADDR => twiddle_h_rsc_0_10_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_10_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_10_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_10_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_10_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_10_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_10_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_10_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_10_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_10_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_10_ARVALID,
      ARREADY => twiddle_h_rsc_0_10_ARREADY,
      RID => twiddle_h_rsc_0_10_i_RID,
      RDATA => twiddle_h_rsc_0_10_i_RDATA,
      RRESP => twiddle_h_rsc_0_10_i_RRESP,
      RLAST => twiddle_h_rsc_0_10_RLAST,
      RUSER => twiddle_h_rsc_0_10_i_RUSER,
      RVALID => twiddle_h_rsc_0_10_RVALID,
      RREADY => twiddle_h_rsc_0_10_RREADY,
      s_re => twiddle_h_rsc_0_10_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_10_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_10_i_s_waddr,
      s_din => twiddle_h_rsc_0_10_i_s_din_1,
      s_dout => twiddle_h_rsc_0_10_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_10_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_10_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_10_is_idle,
      tr_write_done => twiddle_h_rsc_0_10_tr_write_done,
      s_tdone => twiddle_h_rsc_0_10_s_tdone
    );
  twiddle_h_rsc_0_10_i_AWID(0) <= twiddle_h_rsc_0_10_AWID;
  twiddle_h_rsc_0_10_i_AWADDR <= twiddle_h_rsc_0_10_AWADDR;
  twiddle_h_rsc_0_10_i_AWLEN <= twiddle_h_rsc_0_10_AWLEN;
  twiddle_h_rsc_0_10_i_AWSIZE <= twiddle_h_rsc_0_10_AWSIZE;
  twiddle_h_rsc_0_10_i_AWBURST <= twiddle_h_rsc_0_10_AWBURST;
  twiddle_h_rsc_0_10_i_AWCACHE <= twiddle_h_rsc_0_10_AWCACHE;
  twiddle_h_rsc_0_10_i_AWPROT <= twiddle_h_rsc_0_10_AWPROT;
  twiddle_h_rsc_0_10_i_AWQOS <= twiddle_h_rsc_0_10_AWQOS;
  twiddle_h_rsc_0_10_i_AWREGION <= twiddle_h_rsc_0_10_AWREGION;
  twiddle_h_rsc_0_10_i_AWUSER(0) <= twiddle_h_rsc_0_10_AWUSER;
  twiddle_h_rsc_0_10_i_WDATA <= twiddle_h_rsc_0_10_WDATA;
  twiddle_h_rsc_0_10_i_WSTRB <= twiddle_h_rsc_0_10_WSTRB;
  twiddle_h_rsc_0_10_i_WUSER(0) <= twiddle_h_rsc_0_10_WUSER;
  twiddle_h_rsc_0_10_BID <= twiddle_h_rsc_0_10_i_BID(0);
  twiddle_h_rsc_0_10_BRESP <= twiddle_h_rsc_0_10_i_BRESP;
  twiddle_h_rsc_0_10_BUSER <= twiddle_h_rsc_0_10_i_BUSER(0);
  twiddle_h_rsc_0_10_i_ARID(0) <= twiddle_h_rsc_0_10_ARID;
  twiddle_h_rsc_0_10_i_ARADDR <= twiddle_h_rsc_0_10_ARADDR;
  twiddle_h_rsc_0_10_i_ARLEN <= twiddle_h_rsc_0_10_ARLEN;
  twiddle_h_rsc_0_10_i_ARSIZE <= twiddle_h_rsc_0_10_ARSIZE;
  twiddle_h_rsc_0_10_i_ARBURST <= twiddle_h_rsc_0_10_ARBURST;
  twiddle_h_rsc_0_10_i_ARCACHE <= twiddle_h_rsc_0_10_ARCACHE;
  twiddle_h_rsc_0_10_i_ARPROT <= twiddle_h_rsc_0_10_ARPROT;
  twiddle_h_rsc_0_10_i_ARQOS <= twiddle_h_rsc_0_10_ARQOS;
  twiddle_h_rsc_0_10_i_ARREGION <= twiddle_h_rsc_0_10_ARREGION;
  twiddle_h_rsc_0_10_i_ARUSER(0) <= twiddle_h_rsc_0_10_ARUSER;
  twiddle_h_rsc_0_10_RID <= twiddle_h_rsc_0_10_i_RID(0);
  twiddle_h_rsc_0_10_RDATA <= twiddle_h_rsc_0_10_i_RDATA;
  twiddle_h_rsc_0_10_RRESP <= twiddle_h_rsc_0_10_i_RRESP;
  twiddle_h_rsc_0_10_RUSER <= twiddle_h_rsc_0_10_i_RUSER(0);
  twiddle_h_rsc_0_10_i_s_raddr_1 <= twiddle_h_rsc_0_10_i_s_raddr;
  twiddle_h_rsc_0_10_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_10_i_s_din <= twiddle_h_rsc_0_10_i_s_din_1;
  twiddle_h_rsc_0_10_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_10_i_oswt => twiddle_h_rsc_0_10_i_oswt,
      twiddle_h_rsc_0_10_i_biwt => twiddle_h_rsc_0_10_i_biwt,
      twiddle_h_rsc_0_10_i_bdwt => twiddle_h_rsc_0_10_i_bdwt,
      twiddle_h_rsc_0_10_i_bcwt => twiddle_h_rsc_0_10_i_bcwt,
      twiddle_h_rsc_0_10_i_s_re_core_sct => twiddle_h_rsc_0_10_i_s_re_core_sct,
      twiddle_h_rsc_0_10_i_s_rrdy => twiddle_h_rsc_0_10_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_10_i_oswt => twiddle_h_rsc_0_10_i_oswt,
      twiddle_h_rsc_0_10_i_wen_comp => twiddle_h_rsc_0_10_i_wen_comp,
      twiddle_h_rsc_0_10_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp_inst_twiddle_h_rsc_0_10_i_s_raddr_core,
      twiddle_h_rsc_0_10_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp_inst_twiddle_h_rsc_0_10_i_s_din_mxwt,
      twiddle_h_rsc_0_10_i_biwt => twiddle_h_rsc_0_10_i_biwt,
      twiddle_h_rsc_0_10_i_bdwt => twiddle_h_rsc_0_10_i_bdwt,
      twiddle_h_rsc_0_10_i_bcwt => twiddle_h_rsc_0_10_i_bcwt,
      twiddle_h_rsc_0_10_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp_inst_twiddle_h_rsc_0_10_i_s_raddr,
      twiddle_h_rsc_0_10_i_s_raddr_core_sct => twiddle_h_rsc_0_10_i_s_re_core_sct,
      twiddle_h_rsc_0_10_i_s_din => peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp_inst_twiddle_h_rsc_0_10_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp_inst_twiddle_h_rsc_0_10_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_10_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_10_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp_inst_twiddle_h_rsc_0_10_i_s_din_mxwt;
  twiddle_h_rsc_0_10_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp_inst_twiddle_h_rsc_0_10_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_10_i_twiddle_h_rsc_0_10_wait_dp_inst_twiddle_h_rsc_0_10_i_s_din
      <= twiddle_h_rsc_0_10_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_9_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_9_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_9_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_9_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_9_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_9_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_9_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_9_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_9_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_9_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_9_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_9_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_9_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_9_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_9_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_9_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_9_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_9_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_9_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_9_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_9_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_9_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_9_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_9_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_9_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_9_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_9_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_9_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_9_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_9_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_9_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_9_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_9_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_9_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_9_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_9_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_9_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_9_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_9_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_9_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_9_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_9_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_9_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_9_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_9_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_9_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_9_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_9_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_9_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_9_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_9_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_9_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_9_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_9_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_9_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp_inst_twiddle_h_rsc_0_9_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp_inst_twiddle_h_rsc_0_9_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp_inst_twiddle_h_rsc_0_9_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp_inst_twiddle_h_rsc_0_9_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_9_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_9_i_AWID,
      AWADDR => twiddle_h_rsc_0_9_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_9_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_9_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_9_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_9_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_9_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_9_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_9_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_9_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_9_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_9_AWVALID,
      AWREADY => twiddle_h_rsc_0_9_AWREADY,
      WDATA => twiddle_h_rsc_0_9_i_WDATA,
      WSTRB => twiddle_h_rsc_0_9_i_WSTRB,
      WLAST => twiddle_h_rsc_0_9_WLAST,
      WUSER => twiddle_h_rsc_0_9_i_WUSER,
      WVALID => twiddle_h_rsc_0_9_WVALID,
      WREADY => twiddle_h_rsc_0_9_WREADY,
      BID => twiddle_h_rsc_0_9_i_BID,
      BRESP => twiddle_h_rsc_0_9_i_BRESP,
      BUSER => twiddle_h_rsc_0_9_i_BUSER,
      BVALID => twiddle_h_rsc_0_9_BVALID,
      BREADY => twiddle_h_rsc_0_9_BREADY,
      ARID => twiddle_h_rsc_0_9_i_ARID,
      ARADDR => twiddle_h_rsc_0_9_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_9_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_9_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_9_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_9_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_9_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_9_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_9_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_9_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_9_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_9_ARVALID,
      ARREADY => twiddle_h_rsc_0_9_ARREADY,
      RID => twiddle_h_rsc_0_9_i_RID,
      RDATA => twiddle_h_rsc_0_9_i_RDATA,
      RRESP => twiddle_h_rsc_0_9_i_RRESP,
      RLAST => twiddle_h_rsc_0_9_RLAST,
      RUSER => twiddle_h_rsc_0_9_i_RUSER,
      RVALID => twiddle_h_rsc_0_9_RVALID,
      RREADY => twiddle_h_rsc_0_9_RREADY,
      s_re => twiddle_h_rsc_0_9_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_9_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_9_i_s_waddr,
      s_din => twiddle_h_rsc_0_9_i_s_din_1,
      s_dout => twiddle_h_rsc_0_9_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_9_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_9_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_9_is_idle,
      tr_write_done => twiddle_h_rsc_0_9_tr_write_done,
      s_tdone => twiddle_h_rsc_0_9_s_tdone
    );
  twiddle_h_rsc_0_9_i_AWID(0) <= twiddle_h_rsc_0_9_AWID;
  twiddle_h_rsc_0_9_i_AWADDR <= twiddle_h_rsc_0_9_AWADDR;
  twiddle_h_rsc_0_9_i_AWLEN <= twiddle_h_rsc_0_9_AWLEN;
  twiddle_h_rsc_0_9_i_AWSIZE <= twiddle_h_rsc_0_9_AWSIZE;
  twiddle_h_rsc_0_9_i_AWBURST <= twiddle_h_rsc_0_9_AWBURST;
  twiddle_h_rsc_0_9_i_AWCACHE <= twiddle_h_rsc_0_9_AWCACHE;
  twiddle_h_rsc_0_9_i_AWPROT <= twiddle_h_rsc_0_9_AWPROT;
  twiddle_h_rsc_0_9_i_AWQOS <= twiddle_h_rsc_0_9_AWQOS;
  twiddle_h_rsc_0_9_i_AWREGION <= twiddle_h_rsc_0_9_AWREGION;
  twiddle_h_rsc_0_9_i_AWUSER(0) <= twiddle_h_rsc_0_9_AWUSER;
  twiddle_h_rsc_0_9_i_WDATA <= twiddle_h_rsc_0_9_WDATA;
  twiddle_h_rsc_0_9_i_WSTRB <= twiddle_h_rsc_0_9_WSTRB;
  twiddle_h_rsc_0_9_i_WUSER(0) <= twiddle_h_rsc_0_9_WUSER;
  twiddle_h_rsc_0_9_BID <= twiddle_h_rsc_0_9_i_BID(0);
  twiddle_h_rsc_0_9_BRESP <= twiddle_h_rsc_0_9_i_BRESP;
  twiddle_h_rsc_0_9_BUSER <= twiddle_h_rsc_0_9_i_BUSER(0);
  twiddle_h_rsc_0_9_i_ARID(0) <= twiddle_h_rsc_0_9_ARID;
  twiddle_h_rsc_0_9_i_ARADDR <= twiddle_h_rsc_0_9_ARADDR;
  twiddle_h_rsc_0_9_i_ARLEN <= twiddle_h_rsc_0_9_ARLEN;
  twiddle_h_rsc_0_9_i_ARSIZE <= twiddle_h_rsc_0_9_ARSIZE;
  twiddle_h_rsc_0_9_i_ARBURST <= twiddle_h_rsc_0_9_ARBURST;
  twiddle_h_rsc_0_9_i_ARCACHE <= twiddle_h_rsc_0_9_ARCACHE;
  twiddle_h_rsc_0_9_i_ARPROT <= twiddle_h_rsc_0_9_ARPROT;
  twiddle_h_rsc_0_9_i_ARQOS <= twiddle_h_rsc_0_9_ARQOS;
  twiddle_h_rsc_0_9_i_ARREGION <= twiddle_h_rsc_0_9_ARREGION;
  twiddle_h_rsc_0_9_i_ARUSER(0) <= twiddle_h_rsc_0_9_ARUSER;
  twiddle_h_rsc_0_9_RID <= twiddle_h_rsc_0_9_i_RID(0);
  twiddle_h_rsc_0_9_RDATA <= twiddle_h_rsc_0_9_i_RDATA;
  twiddle_h_rsc_0_9_RRESP <= twiddle_h_rsc_0_9_i_RRESP;
  twiddle_h_rsc_0_9_RUSER <= twiddle_h_rsc_0_9_i_RUSER(0);
  twiddle_h_rsc_0_9_i_s_raddr_1 <= twiddle_h_rsc_0_9_i_s_raddr;
  twiddle_h_rsc_0_9_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_9_i_s_din <= twiddle_h_rsc_0_9_i_s_din_1;
  twiddle_h_rsc_0_9_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_9_i_oswt => twiddle_h_rsc_0_9_i_oswt,
      twiddle_h_rsc_0_9_i_biwt => twiddle_h_rsc_0_9_i_biwt,
      twiddle_h_rsc_0_9_i_bdwt => twiddle_h_rsc_0_9_i_bdwt,
      twiddle_h_rsc_0_9_i_bcwt => twiddle_h_rsc_0_9_i_bcwt,
      twiddle_h_rsc_0_9_i_s_re_core_sct => twiddle_h_rsc_0_9_i_s_re_core_sct,
      twiddle_h_rsc_0_9_i_s_rrdy => twiddle_h_rsc_0_9_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_9_i_oswt => twiddle_h_rsc_0_9_i_oswt,
      twiddle_h_rsc_0_9_i_wen_comp => twiddle_h_rsc_0_9_i_wen_comp,
      twiddle_h_rsc_0_9_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp_inst_twiddle_h_rsc_0_9_i_s_raddr_core,
      twiddle_h_rsc_0_9_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp_inst_twiddle_h_rsc_0_9_i_s_din_mxwt,
      twiddle_h_rsc_0_9_i_biwt => twiddle_h_rsc_0_9_i_biwt,
      twiddle_h_rsc_0_9_i_bdwt => twiddle_h_rsc_0_9_i_bdwt,
      twiddle_h_rsc_0_9_i_bcwt => twiddle_h_rsc_0_9_i_bcwt,
      twiddle_h_rsc_0_9_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp_inst_twiddle_h_rsc_0_9_i_s_raddr,
      twiddle_h_rsc_0_9_i_s_raddr_core_sct => twiddle_h_rsc_0_9_i_s_re_core_sct,
      twiddle_h_rsc_0_9_i_s_din => peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp_inst_twiddle_h_rsc_0_9_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp_inst_twiddle_h_rsc_0_9_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_9_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_9_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp_inst_twiddle_h_rsc_0_9_i_s_din_mxwt;
  twiddle_h_rsc_0_9_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp_inst_twiddle_h_rsc_0_9_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_9_i_twiddle_h_rsc_0_9_wait_dp_inst_twiddle_h_rsc_0_9_i_s_din
      <= twiddle_h_rsc_0_9_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_8_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_8_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_8_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_8_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_8_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_8_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_8_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_8_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_8_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_8_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_8_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_8_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_8_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_8_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_8_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_8_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_8_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_8_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_8_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_8_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_8_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_8_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_8_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_8_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_8_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_8_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_8_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_8_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_8_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_8_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_8_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_8_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_8_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_8_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_8_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_8_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_8_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_8_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_8_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_8_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_8_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_8_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_8_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_8_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_8_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_8_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_8_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_8_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_8_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_8_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_8_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_8_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_8_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_8_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_8_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp_inst_twiddle_h_rsc_0_8_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp_inst_twiddle_h_rsc_0_8_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp_inst_twiddle_h_rsc_0_8_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp_inst_twiddle_h_rsc_0_8_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_8_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_8_i_AWID,
      AWADDR => twiddle_h_rsc_0_8_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_8_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_8_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_8_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_8_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_8_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_8_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_8_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_8_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_8_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_8_AWVALID,
      AWREADY => twiddle_h_rsc_0_8_AWREADY,
      WDATA => twiddle_h_rsc_0_8_i_WDATA,
      WSTRB => twiddle_h_rsc_0_8_i_WSTRB,
      WLAST => twiddle_h_rsc_0_8_WLAST,
      WUSER => twiddle_h_rsc_0_8_i_WUSER,
      WVALID => twiddle_h_rsc_0_8_WVALID,
      WREADY => twiddle_h_rsc_0_8_WREADY,
      BID => twiddle_h_rsc_0_8_i_BID,
      BRESP => twiddle_h_rsc_0_8_i_BRESP,
      BUSER => twiddle_h_rsc_0_8_i_BUSER,
      BVALID => twiddle_h_rsc_0_8_BVALID,
      BREADY => twiddle_h_rsc_0_8_BREADY,
      ARID => twiddle_h_rsc_0_8_i_ARID,
      ARADDR => twiddle_h_rsc_0_8_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_8_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_8_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_8_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_8_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_8_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_8_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_8_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_8_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_8_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_8_ARVALID,
      ARREADY => twiddle_h_rsc_0_8_ARREADY,
      RID => twiddle_h_rsc_0_8_i_RID,
      RDATA => twiddle_h_rsc_0_8_i_RDATA,
      RRESP => twiddle_h_rsc_0_8_i_RRESP,
      RLAST => twiddle_h_rsc_0_8_RLAST,
      RUSER => twiddle_h_rsc_0_8_i_RUSER,
      RVALID => twiddle_h_rsc_0_8_RVALID,
      RREADY => twiddle_h_rsc_0_8_RREADY,
      s_re => twiddle_h_rsc_0_8_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_8_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_8_i_s_waddr,
      s_din => twiddle_h_rsc_0_8_i_s_din_1,
      s_dout => twiddle_h_rsc_0_8_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_8_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_8_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_8_is_idle,
      tr_write_done => twiddle_h_rsc_0_8_tr_write_done,
      s_tdone => twiddle_h_rsc_0_8_s_tdone
    );
  twiddle_h_rsc_0_8_i_AWID(0) <= twiddle_h_rsc_0_8_AWID;
  twiddle_h_rsc_0_8_i_AWADDR <= twiddle_h_rsc_0_8_AWADDR;
  twiddle_h_rsc_0_8_i_AWLEN <= twiddle_h_rsc_0_8_AWLEN;
  twiddle_h_rsc_0_8_i_AWSIZE <= twiddle_h_rsc_0_8_AWSIZE;
  twiddle_h_rsc_0_8_i_AWBURST <= twiddle_h_rsc_0_8_AWBURST;
  twiddle_h_rsc_0_8_i_AWCACHE <= twiddle_h_rsc_0_8_AWCACHE;
  twiddle_h_rsc_0_8_i_AWPROT <= twiddle_h_rsc_0_8_AWPROT;
  twiddle_h_rsc_0_8_i_AWQOS <= twiddle_h_rsc_0_8_AWQOS;
  twiddle_h_rsc_0_8_i_AWREGION <= twiddle_h_rsc_0_8_AWREGION;
  twiddle_h_rsc_0_8_i_AWUSER(0) <= twiddle_h_rsc_0_8_AWUSER;
  twiddle_h_rsc_0_8_i_WDATA <= twiddle_h_rsc_0_8_WDATA;
  twiddle_h_rsc_0_8_i_WSTRB <= twiddle_h_rsc_0_8_WSTRB;
  twiddle_h_rsc_0_8_i_WUSER(0) <= twiddle_h_rsc_0_8_WUSER;
  twiddle_h_rsc_0_8_BID <= twiddle_h_rsc_0_8_i_BID(0);
  twiddle_h_rsc_0_8_BRESP <= twiddle_h_rsc_0_8_i_BRESP;
  twiddle_h_rsc_0_8_BUSER <= twiddle_h_rsc_0_8_i_BUSER(0);
  twiddle_h_rsc_0_8_i_ARID(0) <= twiddle_h_rsc_0_8_ARID;
  twiddle_h_rsc_0_8_i_ARADDR <= twiddle_h_rsc_0_8_ARADDR;
  twiddle_h_rsc_0_8_i_ARLEN <= twiddle_h_rsc_0_8_ARLEN;
  twiddle_h_rsc_0_8_i_ARSIZE <= twiddle_h_rsc_0_8_ARSIZE;
  twiddle_h_rsc_0_8_i_ARBURST <= twiddle_h_rsc_0_8_ARBURST;
  twiddle_h_rsc_0_8_i_ARCACHE <= twiddle_h_rsc_0_8_ARCACHE;
  twiddle_h_rsc_0_8_i_ARPROT <= twiddle_h_rsc_0_8_ARPROT;
  twiddle_h_rsc_0_8_i_ARQOS <= twiddle_h_rsc_0_8_ARQOS;
  twiddle_h_rsc_0_8_i_ARREGION <= twiddle_h_rsc_0_8_ARREGION;
  twiddle_h_rsc_0_8_i_ARUSER(0) <= twiddle_h_rsc_0_8_ARUSER;
  twiddle_h_rsc_0_8_RID <= twiddle_h_rsc_0_8_i_RID(0);
  twiddle_h_rsc_0_8_RDATA <= twiddle_h_rsc_0_8_i_RDATA;
  twiddle_h_rsc_0_8_RRESP <= twiddle_h_rsc_0_8_i_RRESP;
  twiddle_h_rsc_0_8_RUSER <= twiddle_h_rsc_0_8_i_RUSER(0);
  twiddle_h_rsc_0_8_i_s_raddr_1 <= twiddle_h_rsc_0_8_i_s_raddr;
  twiddle_h_rsc_0_8_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_8_i_s_din <= twiddle_h_rsc_0_8_i_s_din_1;
  twiddle_h_rsc_0_8_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_8_i_oswt => twiddle_h_rsc_0_8_i_oswt,
      twiddle_h_rsc_0_8_i_biwt => twiddle_h_rsc_0_8_i_biwt,
      twiddle_h_rsc_0_8_i_bdwt => twiddle_h_rsc_0_8_i_bdwt,
      twiddle_h_rsc_0_8_i_bcwt => twiddle_h_rsc_0_8_i_bcwt,
      twiddle_h_rsc_0_8_i_s_re_core_sct => twiddle_h_rsc_0_8_i_s_re_core_sct,
      twiddle_h_rsc_0_8_i_s_rrdy => twiddle_h_rsc_0_8_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_8_i_oswt => twiddle_h_rsc_0_8_i_oswt,
      twiddle_h_rsc_0_8_i_wen_comp => twiddle_h_rsc_0_8_i_wen_comp,
      twiddle_h_rsc_0_8_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp_inst_twiddle_h_rsc_0_8_i_s_raddr_core,
      twiddle_h_rsc_0_8_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp_inst_twiddle_h_rsc_0_8_i_s_din_mxwt,
      twiddle_h_rsc_0_8_i_biwt => twiddle_h_rsc_0_8_i_biwt,
      twiddle_h_rsc_0_8_i_bdwt => twiddle_h_rsc_0_8_i_bdwt,
      twiddle_h_rsc_0_8_i_bcwt => twiddle_h_rsc_0_8_i_bcwt,
      twiddle_h_rsc_0_8_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp_inst_twiddle_h_rsc_0_8_i_s_raddr,
      twiddle_h_rsc_0_8_i_s_raddr_core_sct => twiddle_h_rsc_0_8_i_s_re_core_sct,
      twiddle_h_rsc_0_8_i_s_din => peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp_inst_twiddle_h_rsc_0_8_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp_inst_twiddle_h_rsc_0_8_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_8_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_8_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp_inst_twiddle_h_rsc_0_8_i_s_din_mxwt;
  twiddle_h_rsc_0_8_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp_inst_twiddle_h_rsc_0_8_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_8_i_twiddle_h_rsc_0_8_wait_dp_inst_twiddle_h_rsc_0_8_i_s_din
      <= twiddle_h_rsc_0_8_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_7_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_7_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_7_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_7_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_7_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_7_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_7_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_7_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_7_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_7_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_7_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_7_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_7_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_7_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_7_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_7_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_7_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_7_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_7_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_7_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_7_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_7_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_7_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_7_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_7_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_7_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_7_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_7_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_7_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_7_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_7_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_7_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_7_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_7_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_7_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_7_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_7_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_7_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_7_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_7_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_7_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_7_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_7_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_7_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_7_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_7_i_AWID,
      AWADDR => twiddle_h_rsc_0_7_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_7_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_7_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_7_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_7_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_7_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_7_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_7_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_7_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_7_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_7_AWVALID,
      AWREADY => twiddle_h_rsc_0_7_AWREADY,
      WDATA => twiddle_h_rsc_0_7_i_WDATA,
      WSTRB => twiddle_h_rsc_0_7_i_WSTRB,
      WLAST => twiddle_h_rsc_0_7_WLAST,
      WUSER => twiddle_h_rsc_0_7_i_WUSER,
      WVALID => twiddle_h_rsc_0_7_WVALID,
      WREADY => twiddle_h_rsc_0_7_WREADY,
      BID => twiddle_h_rsc_0_7_i_BID,
      BRESP => twiddle_h_rsc_0_7_i_BRESP,
      BUSER => twiddle_h_rsc_0_7_i_BUSER,
      BVALID => twiddle_h_rsc_0_7_BVALID,
      BREADY => twiddle_h_rsc_0_7_BREADY,
      ARID => twiddle_h_rsc_0_7_i_ARID,
      ARADDR => twiddle_h_rsc_0_7_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_7_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_7_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_7_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_7_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_7_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_7_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_7_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_7_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_7_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_7_ARVALID,
      ARREADY => twiddle_h_rsc_0_7_ARREADY,
      RID => twiddle_h_rsc_0_7_i_RID,
      RDATA => twiddle_h_rsc_0_7_i_RDATA,
      RRESP => twiddle_h_rsc_0_7_i_RRESP,
      RLAST => twiddle_h_rsc_0_7_RLAST,
      RUSER => twiddle_h_rsc_0_7_i_RUSER,
      RVALID => twiddle_h_rsc_0_7_RVALID,
      RREADY => twiddle_h_rsc_0_7_RREADY,
      s_re => twiddle_h_rsc_0_7_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_7_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_7_i_s_waddr,
      s_din => twiddle_h_rsc_0_7_i_s_din_1,
      s_dout => twiddle_h_rsc_0_7_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_7_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_7_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_7_is_idle,
      tr_write_done => twiddle_h_rsc_0_7_tr_write_done,
      s_tdone => twiddle_h_rsc_0_7_s_tdone
    );
  twiddle_h_rsc_0_7_i_AWID(0) <= twiddle_h_rsc_0_7_AWID;
  twiddle_h_rsc_0_7_i_AWADDR <= twiddle_h_rsc_0_7_AWADDR;
  twiddle_h_rsc_0_7_i_AWLEN <= twiddle_h_rsc_0_7_AWLEN;
  twiddle_h_rsc_0_7_i_AWSIZE <= twiddle_h_rsc_0_7_AWSIZE;
  twiddle_h_rsc_0_7_i_AWBURST <= twiddle_h_rsc_0_7_AWBURST;
  twiddle_h_rsc_0_7_i_AWCACHE <= twiddle_h_rsc_0_7_AWCACHE;
  twiddle_h_rsc_0_7_i_AWPROT <= twiddle_h_rsc_0_7_AWPROT;
  twiddle_h_rsc_0_7_i_AWQOS <= twiddle_h_rsc_0_7_AWQOS;
  twiddle_h_rsc_0_7_i_AWREGION <= twiddle_h_rsc_0_7_AWREGION;
  twiddle_h_rsc_0_7_i_AWUSER(0) <= twiddle_h_rsc_0_7_AWUSER;
  twiddle_h_rsc_0_7_i_WDATA <= twiddle_h_rsc_0_7_WDATA;
  twiddle_h_rsc_0_7_i_WSTRB <= twiddle_h_rsc_0_7_WSTRB;
  twiddle_h_rsc_0_7_i_WUSER(0) <= twiddle_h_rsc_0_7_WUSER;
  twiddle_h_rsc_0_7_BID <= twiddle_h_rsc_0_7_i_BID(0);
  twiddle_h_rsc_0_7_BRESP <= twiddle_h_rsc_0_7_i_BRESP;
  twiddle_h_rsc_0_7_BUSER <= twiddle_h_rsc_0_7_i_BUSER(0);
  twiddle_h_rsc_0_7_i_ARID(0) <= twiddle_h_rsc_0_7_ARID;
  twiddle_h_rsc_0_7_i_ARADDR <= twiddle_h_rsc_0_7_ARADDR;
  twiddle_h_rsc_0_7_i_ARLEN <= twiddle_h_rsc_0_7_ARLEN;
  twiddle_h_rsc_0_7_i_ARSIZE <= twiddle_h_rsc_0_7_ARSIZE;
  twiddle_h_rsc_0_7_i_ARBURST <= twiddle_h_rsc_0_7_ARBURST;
  twiddle_h_rsc_0_7_i_ARCACHE <= twiddle_h_rsc_0_7_ARCACHE;
  twiddle_h_rsc_0_7_i_ARPROT <= twiddle_h_rsc_0_7_ARPROT;
  twiddle_h_rsc_0_7_i_ARQOS <= twiddle_h_rsc_0_7_ARQOS;
  twiddle_h_rsc_0_7_i_ARREGION <= twiddle_h_rsc_0_7_ARREGION;
  twiddle_h_rsc_0_7_i_ARUSER(0) <= twiddle_h_rsc_0_7_ARUSER;
  twiddle_h_rsc_0_7_RID <= twiddle_h_rsc_0_7_i_RID(0);
  twiddle_h_rsc_0_7_RDATA <= twiddle_h_rsc_0_7_i_RDATA;
  twiddle_h_rsc_0_7_RRESP <= twiddle_h_rsc_0_7_i_RRESP;
  twiddle_h_rsc_0_7_RUSER <= twiddle_h_rsc_0_7_i_RUSER(0);
  twiddle_h_rsc_0_7_i_s_raddr_1 <= twiddle_h_rsc_0_7_i_s_raddr;
  twiddle_h_rsc_0_7_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_7_i_s_din <= twiddle_h_rsc_0_7_i_s_din_1;
  twiddle_h_rsc_0_7_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_7_i_oswt => twiddle_h_rsc_0_7_i_oswt,
      twiddle_h_rsc_0_7_i_biwt => twiddle_h_rsc_0_7_i_biwt,
      twiddle_h_rsc_0_7_i_bdwt => twiddle_h_rsc_0_7_i_bdwt,
      twiddle_h_rsc_0_7_i_bcwt => twiddle_h_rsc_0_7_i_bcwt,
      twiddle_h_rsc_0_7_i_s_re_core_sct => twiddle_h_rsc_0_7_i_s_re_core_sct,
      twiddle_h_rsc_0_7_i_s_rrdy => twiddle_h_rsc_0_7_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_7_i_oswt => twiddle_h_rsc_0_7_i_oswt,
      twiddle_h_rsc_0_7_i_wen_comp => twiddle_h_rsc_0_7_i_wen_comp,
      twiddle_h_rsc_0_7_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_s_raddr_core,
      twiddle_h_rsc_0_7_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_s_din_mxwt,
      twiddle_h_rsc_0_7_i_biwt => twiddle_h_rsc_0_7_i_biwt,
      twiddle_h_rsc_0_7_i_bdwt => twiddle_h_rsc_0_7_i_bdwt,
      twiddle_h_rsc_0_7_i_bcwt => twiddle_h_rsc_0_7_i_bcwt,
      twiddle_h_rsc_0_7_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_s_raddr,
      twiddle_h_rsc_0_7_i_s_raddr_core_sct => twiddle_h_rsc_0_7_i_s_re_core_sct,
      twiddle_h_rsc_0_7_i_s_din => peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_7_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_7_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_s_din_mxwt;
  twiddle_h_rsc_0_7_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_7_i_twiddle_h_rsc_0_7_wait_dp_inst_twiddle_h_rsc_0_7_i_s_din
      <= twiddle_h_rsc_0_7_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_6_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_6_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_6_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_6_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_6_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_6_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_6_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_6_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_6_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_6_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_6_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_6_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_6_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_6_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_6_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_6_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_6_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_6_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_6_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_6_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_6_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_6_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_6_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_6_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_6_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_6_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_6_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_6_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_6_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_6_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_6_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_6_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_6_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_6_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_6_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_6_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_6_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_6_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_6_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_6_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_6_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_6_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_6_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_6_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_6_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_6_i_AWID,
      AWADDR => twiddle_h_rsc_0_6_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_6_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_6_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_6_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_6_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_6_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_6_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_6_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_6_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_6_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_6_AWVALID,
      AWREADY => twiddle_h_rsc_0_6_AWREADY,
      WDATA => twiddle_h_rsc_0_6_i_WDATA,
      WSTRB => twiddle_h_rsc_0_6_i_WSTRB,
      WLAST => twiddle_h_rsc_0_6_WLAST,
      WUSER => twiddle_h_rsc_0_6_i_WUSER,
      WVALID => twiddle_h_rsc_0_6_WVALID,
      WREADY => twiddle_h_rsc_0_6_WREADY,
      BID => twiddle_h_rsc_0_6_i_BID,
      BRESP => twiddle_h_rsc_0_6_i_BRESP,
      BUSER => twiddle_h_rsc_0_6_i_BUSER,
      BVALID => twiddle_h_rsc_0_6_BVALID,
      BREADY => twiddle_h_rsc_0_6_BREADY,
      ARID => twiddle_h_rsc_0_6_i_ARID,
      ARADDR => twiddle_h_rsc_0_6_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_6_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_6_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_6_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_6_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_6_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_6_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_6_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_6_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_6_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_6_ARVALID,
      ARREADY => twiddle_h_rsc_0_6_ARREADY,
      RID => twiddle_h_rsc_0_6_i_RID,
      RDATA => twiddle_h_rsc_0_6_i_RDATA,
      RRESP => twiddle_h_rsc_0_6_i_RRESP,
      RLAST => twiddle_h_rsc_0_6_RLAST,
      RUSER => twiddle_h_rsc_0_6_i_RUSER,
      RVALID => twiddle_h_rsc_0_6_RVALID,
      RREADY => twiddle_h_rsc_0_6_RREADY,
      s_re => twiddle_h_rsc_0_6_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_6_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_6_i_s_waddr,
      s_din => twiddle_h_rsc_0_6_i_s_din_1,
      s_dout => twiddle_h_rsc_0_6_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_6_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_6_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_6_is_idle,
      tr_write_done => twiddle_h_rsc_0_6_tr_write_done,
      s_tdone => twiddle_h_rsc_0_6_s_tdone
    );
  twiddle_h_rsc_0_6_i_AWID(0) <= twiddle_h_rsc_0_6_AWID;
  twiddle_h_rsc_0_6_i_AWADDR <= twiddle_h_rsc_0_6_AWADDR;
  twiddle_h_rsc_0_6_i_AWLEN <= twiddle_h_rsc_0_6_AWLEN;
  twiddle_h_rsc_0_6_i_AWSIZE <= twiddle_h_rsc_0_6_AWSIZE;
  twiddle_h_rsc_0_6_i_AWBURST <= twiddle_h_rsc_0_6_AWBURST;
  twiddle_h_rsc_0_6_i_AWCACHE <= twiddle_h_rsc_0_6_AWCACHE;
  twiddle_h_rsc_0_6_i_AWPROT <= twiddle_h_rsc_0_6_AWPROT;
  twiddle_h_rsc_0_6_i_AWQOS <= twiddle_h_rsc_0_6_AWQOS;
  twiddle_h_rsc_0_6_i_AWREGION <= twiddle_h_rsc_0_6_AWREGION;
  twiddle_h_rsc_0_6_i_AWUSER(0) <= twiddle_h_rsc_0_6_AWUSER;
  twiddle_h_rsc_0_6_i_WDATA <= twiddle_h_rsc_0_6_WDATA;
  twiddle_h_rsc_0_6_i_WSTRB <= twiddle_h_rsc_0_6_WSTRB;
  twiddle_h_rsc_0_6_i_WUSER(0) <= twiddle_h_rsc_0_6_WUSER;
  twiddle_h_rsc_0_6_BID <= twiddle_h_rsc_0_6_i_BID(0);
  twiddle_h_rsc_0_6_BRESP <= twiddle_h_rsc_0_6_i_BRESP;
  twiddle_h_rsc_0_6_BUSER <= twiddle_h_rsc_0_6_i_BUSER(0);
  twiddle_h_rsc_0_6_i_ARID(0) <= twiddle_h_rsc_0_6_ARID;
  twiddle_h_rsc_0_6_i_ARADDR <= twiddle_h_rsc_0_6_ARADDR;
  twiddle_h_rsc_0_6_i_ARLEN <= twiddle_h_rsc_0_6_ARLEN;
  twiddle_h_rsc_0_6_i_ARSIZE <= twiddle_h_rsc_0_6_ARSIZE;
  twiddle_h_rsc_0_6_i_ARBURST <= twiddle_h_rsc_0_6_ARBURST;
  twiddle_h_rsc_0_6_i_ARCACHE <= twiddle_h_rsc_0_6_ARCACHE;
  twiddle_h_rsc_0_6_i_ARPROT <= twiddle_h_rsc_0_6_ARPROT;
  twiddle_h_rsc_0_6_i_ARQOS <= twiddle_h_rsc_0_6_ARQOS;
  twiddle_h_rsc_0_6_i_ARREGION <= twiddle_h_rsc_0_6_ARREGION;
  twiddle_h_rsc_0_6_i_ARUSER(0) <= twiddle_h_rsc_0_6_ARUSER;
  twiddle_h_rsc_0_6_RID <= twiddle_h_rsc_0_6_i_RID(0);
  twiddle_h_rsc_0_6_RDATA <= twiddle_h_rsc_0_6_i_RDATA;
  twiddle_h_rsc_0_6_RRESP <= twiddle_h_rsc_0_6_i_RRESP;
  twiddle_h_rsc_0_6_RUSER <= twiddle_h_rsc_0_6_i_RUSER(0);
  twiddle_h_rsc_0_6_i_s_raddr_1 <= twiddle_h_rsc_0_6_i_s_raddr;
  twiddle_h_rsc_0_6_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_6_i_s_din <= twiddle_h_rsc_0_6_i_s_din_1;
  twiddle_h_rsc_0_6_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_6_i_oswt => twiddle_h_rsc_0_6_i_oswt,
      twiddle_h_rsc_0_6_i_biwt => twiddle_h_rsc_0_6_i_biwt,
      twiddle_h_rsc_0_6_i_bdwt => twiddle_h_rsc_0_6_i_bdwt,
      twiddle_h_rsc_0_6_i_bcwt => twiddle_h_rsc_0_6_i_bcwt,
      twiddle_h_rsc_0_6_i_s_re_core_sct => twiddle_h_rsc_0_6_i_s_re_core_sct,
      twiddle_h_rsc_0_6_i_s_rrdy => twiddle_h_rsc_0_6_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_6_i_oswt => twiddle_h_rsc_0_6_i_oswt,
      twiddle_h_rsc_0_6_i_wen_comp => twiddle_h_rsc_0_6_i_wen_comp,
      twiddle_h_rsc_0_6_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_s_raddr_core,
      twiddle_h_rsc_0_6_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_s_din_mxwt,
      twiddle_h_rsc_0_6_i_biwt => twiddle_h_rsc_0_6_i_biwt,
      twiddle_h_rsc_0_6_i_bdwt => twiddle_h_rsc_0_6_i_bdwt,
      twiddle_h_rsc_0_6_i_bcwt => twiddle_h_rsc_0_6_i_bcwt,
      twiddle_h_rsc_0_6_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_s_raddr,
      twiddle_h_rsc_0_6_i_s_raddr_core_sct => twiddle_h_rsc_0_6_i_s_re_core_sct,
      twiddle_h_rsc_0_6_i_s_din => peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_6_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_6_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_s_din_mxwt;
  twiddle_h_rsc_0_6_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_6_i_twiddle_h_rsc_0_6_wait_dp_inst_twiddle_h_rsc_0_6_i_s_din
      <= twiddle_h_rsc_0_6_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_5_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_5_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_5_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_5_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_5_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_5_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_5_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_5_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_5_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_5_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_5_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_5_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_5_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_5_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_5_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_5_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_5_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_5_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_5_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_5_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_5_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_5_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_5_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_5_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_5_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_5_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_5_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_5_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_5_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_5_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_5_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_5_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_5_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_5_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_5_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_5_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_5_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_5_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_5_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_5_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_5_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_5_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_5_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_5_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_5_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_5_i_AWID,
      AWADDR => twiddle_h_rsc_0_5_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_5_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_5_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_5_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_5_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_5_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_5_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_5_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_5_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_5_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_5_AWVALID,
      AWREADY => twiddle_h_rsc_0_5_AWREADY,
      WDATA => twiddle_h_rsc_0_5_i_WDATA,
      WSTRB => twiddle_h_rsc_0_5_i_WSTRB,
      WLAST => twiddle_h_rsc_0_5_WLAST,
      WUSER => twiddle_h_rsc_0_5_i_WUSER,
      WVALID => twiddle_h_rsc_0_5_WVALID,
      WREADY => twiddle_h_rsc_0_5_WREADY,
      BID => twiddle_h_rsc_0_5_i_BID,
      BRESP => twiddle_h_rsc_0_5_i_BRESP,
      BUSER => twiddle_h_rsc_0_5_i_BUSER,
      BVALID => twiddle_h_rsc_0_5_BVALID,
      BREADY => twiddle_h_rsc_0_5_BREADY,
      ARID => twiddle_h_rsc_0_5_i_ARID,
      ARADDR => twiddle_h_rsc_0_5_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_5_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_5_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_5_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_5_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_5_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_5_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_5_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_5_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_5_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_5_ARVALID,
      ARREADY => twiddle_h_rsc_0_5_ARREADY,
      RID => twiddle_h_rsc_0_5_i_RID,
      RDATA => twiddle_h_rsc_0_5_i_RDATA,
      RRESP => twiddle_h_rsc_0_5_i_RRESP,
      RLAST => twiddle_h_rsc_0_5_RLAST,
      RUSER => twiddle_h_rsc_0_5_i_RUSER,
      RVALID => twiddle_h_rsc_0_5_RVALID,
      RREADY => twiddle_h_rsc_0_5_RREADY,
      s_re => twiddle_h_rsc_0_5_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_5_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_5_i_s_waddr,
      s_din => twiddle_h_rsc_0_5_i_s_din_1,
      s_dout => twiddle_h_rsc_0_5_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_5_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_5_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_5_is_idle,
      tr_write_done => twiddle_h_rsc_0_5_tr_write_done,
      s_tdone => twiddle_h_rsc_0_5_s_tdone
    );
  twiddle_h_rsc_0_5_i_AWID(0) <= twiddle_h_rsc_0_5_AWID;
  twiddle_h_rsc_0_5_i_AWADDR <= twiddle_h_rsc_0_5_AWADDR;
  twiddle_h_rsc_0_5_i_AWLEN <= twiddle_h_rsc_0_5_AWLEN;
  twiddle_h_rsc_0_5_i_AWSIZE <= twiddle_h_rsc_0_5_AWSIZE;
  twiddle_h_rsc_0_5_i_AWBURST <= twiddle_h_rsc_0_5_AWBURST;
  twiddle_h_rsc_0_5_i_AWCACHE <= twiddle_h_rsc_0_5_AWCACHE;
  twiddle_h_rsc_0_5_i_AWPROT <= twiddle_h_rsc_0_5_AWPROT;
  twiddle_h_rsc_0_5_i_AWQOS <= twiddle_h_rsc_0_5_AWQOS;
  twiddle_h_rsc_0_5_i_AWREGION <= twiddle_h_rsc_0_5_AWREGION;
  twiddle_h_rsc_0_5_i_AWUSER(0) <= twiddle_h_rsc_0_5_AWUSER;
  twiddle_h_rsc_0_5_i_WDATA <= twiddle_h_rsc_0_5_WDATA;
  twiddle_h_rsc_0_5_i_WSTRB <= twiddle_h_rsc_0_5_WSTRB;
  twiddle_h_rsc_0_5_i_WUSER(0) <= twiddle_h_rsc_0_5_WUSER;
  twiddle_h_rsc_0_5_BID <= twiddle_h_rsc_0_5_i_BID(0);
  twiddle_h_rsc_0_5_BRESP <= twiddle_h_rsc_0_5_i_BRESP;
  twiddle_h_rsc_0_5_BUSER <= twiddle_h_rsc_0_5_i_BUSER(0);
  twiddle_h_rsc_0_5_i_ARID(0) <= twiddle_h_rsc_0_5_ARID;
  twiddle_h_rsc_0_5_i_ARADDR <= twiddle_h_rsc_0_5_ARADDR;
  twiddle_h_rsc_0_5_i_ARLEN <= twiddle_h_rsc_0_5_ARLEN;
  twiddle_h_rsc_0_5_i_ARSIZE <= twiddle_h_rsc_0_5_ARSIZE;
  twiddle_h_rsc_0_5_i_ARBURST <= twiddle_h_rsc_0_5_ARBURST;
  twiddle_h_rsc_0_5_i_ARCACHE <= twiddle_h_rsc_0_5_ARCACHE;
  twiddle_h_rsc_0_5_i_ARPROT <= twiddle_h_rsc_0_5_ARPROT;
  twiddle_h_rsc_0_5_i_ARQOS <= twiddle_h_rsc_0_5_ARQOS;
  twiddle_h_rsc_0_5_i_ARREGION <= twiddle_h_rsc_0_5_ARREGION;
  twiddle_h_rsc_0_5_i_ARUSER(0) <= twiddle_h_rsc_0_5_ARUSER;
  twiddle_h_rsc_0_5_RID <= twiddle_h_rsc_0_5_i_RID(0);
  twiddle_h_rsc_0_5_RDATA <= twiddle_h_rsc_0_5_i_RDATA;
  twiddle_h_rsc_0_5_RRESP <= twiddle_h_rsc_0_5_i_RRESP;
  twiddle_h_rsc_0_5_RUSER <= twiddle_h_rsc_0_5_i_RUSER(0);
  twiddle_h_rsc_0_5_i_s_raddr_1 <= twiddle_h_rsc_0_5_i_s_raddr;
  twiddle_h_rsc_0_5_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_5_i_s_din <= twiddle_h_rsc_0_5_i_s_din_1;
  twiddle_h_rsc_0_5_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_5_i_oswt => twiddle_h_rsc_0_5_i_oswt,
      twiddle_h_rsc_0_5_i_biwt => twiddle_h_rsc_0_5_i_biwt,
      twiddle_h_rsc_0_5_i_bdwt => twiddle_h_rsc_0_5_i_bdwt,
      twiddle_h_rsc_0_5_i_bcwt => twiddle_h_rsc_0_5_i_bcwt,
      twiddle_h_rsc_0_5_i_s_re_core_sct => twiddle_h_rsc_0_5_i_s_re_core_sct,
      twiddle_h_rsc_0_5_i_s_rrdy => twiddle_h_rsc_0_5_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_5_i_oswt => twiddle_h_rsc_0_5_i_oswt,
      twiddle_h_rsc_0_5_i_wen_comp => twiddle_h_rsc_0_5_i_wen_comp,
      twiddle_h_rsc_0_5_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_s_raddr_core,
      twiddle_h_rsc_0_5_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_s_din_mxwt,
      twiddle_h_rsc_0_5_i_biwt => twiddle_h_rsc_0_5_i_biwt,
      twiddle_h_rsc_0_5_i_bdwt => twiddle_h_rsc_0_5_i_bdwt,
      twiddle_h_rsc_0_5_i_bcwt => twiddle_h_rsc_0_5_i_bcwt,
      twiddle_h_rsc_0_5_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_s_raddr,
      twiddle_h_rsc_0_5_i_s_raddr_core_sct => twiddle_h_rsc_0_5_i_s_re_core_sct,
      twiddle_h_rsc_0_5_i_s_din => peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_5_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_5_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_s_din_mxwt;
  twiddle_h_rsc_0_5_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_5_i_twiddle_h_rsc_0_5_wait_dp_inst_twiddle_h_rsc_0_5_i_s_din
      <= twiddle_h_rsc_0_5_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_4_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_4_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_4_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_4_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_4_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_4_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_4_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_4_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_4_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_4_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_4_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_4_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_4_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_4_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_4_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_4_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_4_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_4_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_4_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_4_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_4_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_4_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_4_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_4_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_4_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_4_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_4_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_4_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_4_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_4_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_4_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_4_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_4_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_4_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_4_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_4_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_4_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_4_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_4_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_4_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_4_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_4_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_4_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_4_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_4_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_4_i_AWID,
      AWADDR => twiddle_h_rsc_0_4_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_4_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_4_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_4_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_4_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_4_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_4_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_4_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_4_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_4_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_4_AWVALID,
      AWREADY => twiddle_h_rsc_0_4_AWREADY,
      WDATA => twiddle_h_rsc_0_4_i_WDATA,
      WSTRB => twiddle_h_rsc_0_4_i_WSTRB,
      WLAST => twiddle_h_rsc_0_4_WLAST,
      WUSER => twiddle_h_rsc_0_4_i_WUSER,
      WVALID => twiddle_h_rsc_0_4_WVALID,
      WREADY => twiddle_h_rsc_0_4_WREADY,
      BID => twiddle_h_rsc_0_4_i_BID,
      BRESP => twiddle_h_rsc_0_4_i_BRESP,
      BUSER => twiddle_h_rsc_0_4_i_BUSER,
      BVALID => twiddle_h_rsc_0_4_BVALID,
      BREADY => twiddle_h_rsc_0_4_BREADY,
      ARID => twiddle_h_rsc_0_4_i_ARID,
      ARADDR => twiddle_h_rsc_0_4_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_4_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_4_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_4_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_4_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_4_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_4_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_4_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_4_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_4_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_4_ARVALID,
      ARREADY => twiddle_h_rsc_0_4_ARREADY,
      RID => twiddle_h_rsc_0_4_i_RID,
      RDATA => twiddle_h_rsc_0_4_i_RDATA,
      RRESP => twiddle_h_rsc_0_4_i_RRESP,
      RLAST => twiddle_h_rsc_0_4_RLAST,
      RUSER => twiddle_h_rsc_0_4_i_RUSER,
      RVALID => twiddle_h_rsc_0_4_RVALID,
      RREADY => twiddle_h_rsc_0_4_RREADY,
      s_re => twiddle_h_rsc_0_4_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_4_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_4_i_s_waddr,
      s_din => twiddle_h_rsc_0_4_i_s_din_1,
      s_dout => twiddle_h_rsc_0_4_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_4_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_4_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_4_is_idle,
      tr_write_done => twiddle_h_rsc_0_4_tr_write_done,
      s_tdone => twiddle_h_rsc_0_4_s_tdone
    );
  twiddle_h_rsc_0_4_i_AWID(0) <= twiddle_h_rsc_0_4_AWID;
  twiddle_h_rsc_0_4_i_AWADDR <= twiddle_h_rsc_0_4_AWADDR;
  twiddle_h_rsc_0_4_i_AWLEN <= twiddle_h_rsc_0_4_AWLEN;
  twiddle_h_rsc_0_4_i_AWSIZE <= twiddle_h_rsc_0_4_AWSIZE;
  twiddle_h_rsc_0_4_i_AWBURST <= twiddle_h_rsc_0_4_AWBURST;
  twiddle_h_rsc_0_4_i_AWCACHE <= twiddle_h_rsc_0_4_AWCACHE;
  twiddle_h_rsc_0_4_i_AWPROT <= twiddle_h_rsc_0_4_AWPROT;
  twiddle_h_rsc_0_4_i_AWQOS <= twiddle_h_rsc_0_4_AWQOS;
  twiddle_h_rsc_0_4_i_AWREGION <= twiddle_h_rsc_0_4_AWREGION;
  twiddle_h_rsc_0_4_i_AWUSER(0) <= twiddle_h_rsc_0_4_AWUSER;
  twiddle_h_rsc_0_4_i_WDATA <= twiddle_h_rsc_0_4_WDATA;
  twiddle_h_rsc_0_4_i_WSTRB <= twiddle_h_rsc_0_4_WSTRB;
  twiddle_h_rsc_0_4_i_WUSER(0) <= twiddle_h_rsc_0_4_WUSER;
  twiddle_h_rsc_0_4_BID <= twiddle_h_rsc_0_4_i_BID(0);
  twiddle_h_rsc_0_4_BRESP <= twiddle_h_rsc_0_4_i_BRESP;
  twiddle_h_rsc_0_4_BUSER <= twiddle_h_rsc_0_4_i_BUSER(0);
  twiddle_h_rsc_0_4_i_ARID(0) <= twiddle_h_rsc_0_4_ARID;
  twiddle_h_rsc_0_4_i_ARADDR <= twiddle_h_rsc_0_4_ARADDR;
  twiddle_h_rsc_0_4_i_ARLEN <= twiddle_h_rsc_0_4_ARLEN;
  twiddle_h_rsc_0_4_i_ARSIZE <= twiddle_h_rsc_0_4_ARSIZE;
  twiddle_h_rsc_0_4_i_ARBURST <= twiddle_h_rsc_0_4_ARBURST;
  twiddle_h_rsc_0_4_i_ARCACHE <= twiddle_h_rsc_0_4_ARCACHE;
  twiddle_h_rsc_0_4_i_ARPROT <= twiddle_h_rsc_0_4_ARPROT;
  twiddle_h_rsc_0_4_i_ARQOS <= twiddle_h_rsc_0_4_ARQOS;
  twiddle_h_rsc_0_4_i_ARREGION <= twiddle_h_rsc_0_4_ARREGION;
  twiddle_h_rsc_0_4_i_ARUSER(0) <= twiddle_h_rsc_0_4_ARUSER;
  twiddle_h_rsc_0_4_RID <= twiddle_h_rsc_0_4_i_RID(0);
  twiddle_h_rsc_0_4_RDATA <= twiddle_h_rsc_0_4_i_RDATA;
  twiddle_h_rsc_0_4_RRESP <= twiddle_h_rsc_0_4_i_RRESP;
  twiddle_h_rsc_0_4_RUSER <= twiddle_h_rsc_0_4_i_RUSER(0);
  twiddle_h_rsc_0_4_i_s_raddr_1 <= twiddle_h_rsc_0_4_i_s_raddr;
  twiddle_h_rsc_0_4_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_4_i_s_din <= twiddle_h_rsc_0_4_i_s_din_1;
  twiddle_h_rsc_0_4_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_4_i_oswt => twiddle_h_rsc_0_4_i_oswt,
      twiddle_h_rsc_0_4_i_biwt => twiddle_h_rsc_0_4_i_biwt,
      twiddle_h_rsc_0_4_i_bdwt => twiddle_h_rsc_0_4_i_bdwt,
      twiddle_h_rsc_0_4_i_bcwt => twiddle_h_rsc_0_4_i_bcwt,
      twiddle_h_rsc_0_4_i_s_re_core_sct => twiddle_h_rsc_0_4_i_s_re_core_sct,
      twiddle_h_rsc_0_4_i_s_rrdy => twiddle_h_rsc_0_4_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_4_i_oswt => twiddle_h_rsc_0_4_i_oswt,
      twiddle_h_rsc_0_4_i_wen_comp => twiddle_h_rsc_0_4_i_wen_comp,
      twiddle_h_rsc_0_4_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_s_raddr_core,
      twiddle_h_rsc_0_4_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_s_din_mxwt,
      twiddle_h_rsc_0_4_i_biwt => twiddle_h_rsc_0_4_i_biwt,
      twiddle_h_rsc_0_4_i_bdwt => twiddle_h_rsc_0_4_i_bdwt,
      twiddle_h_rsc_0_4_i_bcwt => twiddle_h_rsc_0_4_i_bcwt,
      twiddle_h_rsc_0_4_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_s_raddr,
      twiddle_h_rsc_0_4_i_s_raddr_core_sct => twiddle_h_rsc_0_4_i_s_re_core_sct,
      twiddle_h_rsc_0_4_i_s_din => peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_4_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_4_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_s_din_mxwt;
  twiddle_h_rsc_0_4_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_4_i_twiddle_h_rsc_0_4_wait_dp_inst_twiddle_h_rsc_0_4_i_s_din
      <= twiddle_h_rsc_0_4_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_3_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_3_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_3_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_3_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_3_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_3_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_3_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_3_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_3_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_3_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_3_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_3_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_3_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_3_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_3_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_3_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_3_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_3_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_3_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_3_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_3_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_3_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_3_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_3_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_3_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_3_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_3_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_3_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_3_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_3_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_3_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_3_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_3_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_3_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_3_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_3_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_3_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_3_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_3_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_3_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_3_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_3_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_3_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_3_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_3_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_3_i_AWID,
      AWADDR => twiddle_h_rsc_0_3_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_3_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_3_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_3_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_3_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_3_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_3_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_3_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_3_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_3_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_3_AWVALID,
      AWREADY => twiddle_h_rsc_0_3_AWREADY,
      WDATA => twiddle_h_rsc_0_3_i_WDATA,
      WSTRB => twiddle_h_rsc_0_3_i_WSTRB,
      WLAST => twiddle_h_rsc_0_3_WLAST,
      WUSER => twiddle_h_rsc_0_3_i_WUSER,
      WVALID => twiddle_h_rsc_0_3_WVALID,
      WREADY => twiddle_h_rsc_0_3_WREADY,
      BID => twiddle_h_rsc_0_3_i_BID,
      BRESP => twiddle_h_rsc_0_3_i_BRESP,
      BUSER => twiddle_h_rsc_0_3_i_BUSER,
      BVALID => twiddle_h_rsc_0_3_BVALID,
      BREADY => twiddle_h_rsc_0_3_BREADY,
      ARID => twiddle_h_rsc_0_3_i_ARID,
      ARADDR => twiddle_h_rsc_0_3_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_3_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_3_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_3_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_3_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_3_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_3_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_3_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_3_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_3_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_3_ARVALID,
      ARREADY => twiddle_h_rsc_0_3_ARREADY,
      RID => twiddle_h_rsc_0_3_i_RID,
      RDATA => twiddle_h_rsc_0_3_i_RDATA,
      RRESP => twiddle_h_rsc_0_3_i_RRESP,
      RLAST => twiddle_h_rsc_0_3_RLAST,
      RUSER => twiddle_h_rsc_0_3_i_RUSER,
      RVALID => twiddle_h_rsc_0_3_RVALID,
      RREADY => twiddle_h_rsc_0_3_RREADY,
      s_re => twiddle_h_rsc_0_3_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_3_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_3_i_s_waddr,
      s_din => twiddle_h_rsc_0_3_i_s_din_1,
      s_dout => twiddle_h_rsc_0_3_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_3_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_3_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_3_is_idle,
      tr_write_done => twiddle_h_rsc_0_3_tr_write_done,
      s_tdone => twiddle_h_rsc_0_3_s_tdone
    );
  twiddle_h_rsc_0_3_i_AWID(0) <= twiddle_h_rsc_0_3_AWID;
  twiddle_h_rsc_0_3_i_AWADDR <= twiddle_h_rsc_0_3_AWADDR;
  twiddle_h_rsc_0_3_i_AWLEN <= twiddle_h_rsc_0_3_AWLEN;
  twiddle_h_rsc_0_3_i_AWSIZE <= twiddle_h_rsc_0_3_AWSIZE;
  twiddle_h_rsc_0_3_i_AWBURST <= twiddle_h_rsc_0_3_AWBURST;
  twiddle_h_rsc_0_3_i_AWCACHE <= twiddle_h_rsc_0_3_AWCACHE;
  twiddle_h_rsc_0_3_i_AWPROT <= twiddle_h_rsc_0_3_AWPROT;
  twiddle_h_rsc_0_3_i_AWQOS <= twiddle_h_rsc_0_3_AWQOS;
  twiddle_h_rsc_0_3_i_AWREGION <= twiddle_h_rsc_0_3_AWREGION;
  twiddle_h_rsc_0_3_i_AWUSER(0) <= twiddle_h_rsc_0_3_AWUSER;
  twiddle_h_rsc_0_3_i_WDATA <= twiddle_h_rsc_0_3_WDATA;
  twiddle_h_rsc_0_3_i_WSTRB <= twiddle_h_rsc_0_3_WSTRB;
  twiddle_h_rsc_0_3_i_WUSER(0) <= twiddle_h_rsc_0_3_WUSER;
  twiddle_h_rsc_0_3_BID <= twiddle_h_rsc_0_3_i_BID(0);
  twiddle_h_rsc_0_3_BRESP <= twiddle_h_rsc_0_3_i_BRESP;
  twiddle_h_rsc_0_3_BUSER <= twiddle_h_rsc_0_3_i_BUSER(0);
  twiddle_h_rsc_0_3_i_ARID(0) <= twiddle_h_rsc_0_3_ARID;
  twiddle_h_rsc_0_3_i_ARADDR <= twiddle_h_rsc_0_3_ARADDR;
  twiddle_h_rsc_0_3_i_ARLEN <= twiddle_h_rsc_0_3_ARLEN;
  twiddle_h_rsc_0_3_i_ARSIZE <= twiddle_h_rsc_0_3_ARSIZE;
  twiddle_h_rsc_0_3_i_ARBURST <= twiddle_h_rsc_0_3_ARBURST;
  twiddle_h_rsc_0_3_i_ARCACHE <= twiddle_h_rsc_0_3_ARCACHE;
  twiddle_h_rsc_0_3_i_ARPROT <= twiddle_h_rsc_0_3_ARPROT;
  twiddle_h_rsc_0_3_i_ARQOS <= twiddle_h_rsc_0_3_ARQOS;
  twiddle_h_rsc_0_3_i_ARREGION <= twiddle_h_rsc_0_3_ARREGION;
  twiddle_h_rsc_0_3_i_ARUSER(0) <= twiddle_h_rsc_0_3_ARUSER;
  twiddle_h_rsc_0_3_RID <= twiddle_h_rsc_0_3_i_RID(0);
  twiddle_h_rsc_0_3_RDATA <= twiddle_h_rsc_0_3_i_RDATA;
  twiddle_h_rsc_0_3_RRESP <= twiddle_h_rsc_0_3_i_RRESP;
  twiddle_h_rsc_0_3_RUSER <= twiddle_h_rsc_0_3_i_RUSER(0);
  twiddle_h_rsc_0_3_i_s_raddr_1 <= twiddle_h_rsc_0_3_i_s_raddr;
  twiddle_h_rsc_0_3_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_3_i_s_din <= twiddle_h_rsc_0_3_i_s_din_1;
  twiddle_h_rsc_0_3_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_3_i_oswt => twiddle_h_rsc_0_3_i_oswt,
      twiddle_h_rsc_0_3_i_biwt => twiddle_h_rsc_0_3_i_biwt,
      twiddle_h_rsc_0_3_i_bdwt => twiddle_h_rsc_0_3_i_bdwt,
      twiddle_h_rsc_0_3_i_bcwt => twiddle_h_rsc_0_3_i_bcwt,
      twiddle_h_rsc_0_3_i_s_re_core_sct => twiddle_h_rsc_0_3_i_s_re_core_sct,
      twiddle_h_rsc_0_3_i_s_rrdy => twiddle_h_rsc_0_3_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_3_i_oswt => twiddle_h_rsc_0_3_i_oswt,
      twiddle_h_rsc_0_3_i_wen_comp => twiddle_h_rsc_0_3_i_wen_comp,
      twiddle_h_rsc_0_3_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_s_raddr_core,
      twiddle_h_rsc_0_3_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_s_din_mxwt,
      twiddle_h_rsc_0_3_i_biwt => twiddle_h_rsc_0_3_i_biwt,
      twiddle_h_rsc_0_3_i_bdwt => twiddle_h_rsc_0_3_i_bdwt,
      twiddle_h_rsc_0_3_i_bcwt => twiddle_h_rsc_0_3_i_bcwt,
      twiddle_h_rsc_0_3_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_s_raddr,
      twiddle_h_rsc_0_3_i_s_raddr_core_sct => twiddle_h_rsc_0_3_i_s_re_core_sct,
      twiddle_h_rsc_0_3_i_s_din => peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_3_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_3_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_s_din_mxwt;
  twiddle_h_rsc_0_3_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_3_i_twiddle_h_rsc_0_3_wait_dp_inst_twiddle_h_rsc_0_3_i_s_din
      <= twiddle_h_rsc_0_3_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_2_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_2_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_2_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_2_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_2_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_2_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_2_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_2_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_2_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_2_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_2_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_2_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_2_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_2_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_2_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_2_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_2_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_2_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_2_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_2_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_2_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_2_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_2_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_2_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_2_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_2_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_2_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_2_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_2_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_2_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_2_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_2_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_2_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_2_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_2_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_2_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_2_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_2_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_2_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_2_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_2_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_2_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_2_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_2_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_2_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_2_i_AWID,
      AWADDR => twiddle_h_rsc_0_2_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_2_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_2_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_2_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_2_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_2_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_2_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_2_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_2_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_2_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_2_AWVALID,
      AWREADY => twiddle_h_rsc_0_2_AWREADY,
      WDATA => twiddle_h_rsc_0_2_i_WDATA,
      WSTRB => twiddle_h_rsc_0_2_i_WSTRB,
      WLAST => twiddle_h_rsc_0_2_WLAST,
      WUSER => twiddle_h_rsc_0_2_i_WUSER,
      WVALID => twiddle_h_rsc_0_2_WVALID,
      WREADY => twiddle_h_rsc_0_2_WREADY,
      BID => twiddle_h_rsc_0_2_i_BID,
      BRESP => twiddle_h_rsc_0_2_i_BRESP,
      BUSER => twiddle_h_rsc_0_2_i_BUSER,
      BVALID => twiddle_h_rsc_0_2_BVALID,
      BREADY => twiddle_h_rsc_0_2_BREADY,
      ARID => twiddle_h_rsc_0_2_i_ARID,
      ARADDR => twiddle_h_rsc_0_2_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_2_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_2_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_2_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_2_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_2_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_2_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_2_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_2_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_2_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_2_ARVALID,
      ARREADY => twiddle_h_rsc_0_2_ARREADY,
      RID => twiddle_h_rsc_0_2_i_RID,
      RDATA => twiddle_h_rsc_0_2_i_RDATA,
      RRESP => twiddle_h_rsc_0_2_i_RRESP,
      RLAST => twiddle_h_rsc_0_2_RLAST,
      RUSER => twiddle_h_rsc_0_2_i_RUSER,
      RVALID => twiddle_h_rsc_0_2_RVALID,
      RREADY => twiddle_h_rsc_0_2_RREADY,
      s_re => twiddle_h_rsc_0_2_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_2_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_2_i_s_waddr,
      s_din => twiddle_h_rsc_0_2_i_s_din_1,
      s_dout => twiddle_h_rsc_0_2_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_2_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_2_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_2_is_idle,
      tr_write_done => twiddle_h_rsc_0_2_tr_write_done,
      s_tdone => twiddle_h_rsc_0_2_s_tdone
    );
  twiddle_h_rsc_0_2_i_AWID(0) <= twiddle_h_rsc_0_2_AWID;
  twiddle_h_rsc_0_2_i_AWADDR <= twiddle_h_rsc_0_2_AWADDR;
  twiddle_h_rsc_0_2_i_AWLEN <= twiddle_h_rsc_0_2_AWLEN;
  twiddle_h_rsc_0_2_i_AWSIZE <= twiddle_h_rsc_0_2_AWSIZE;
  twiddle_h_rsc_0_2_i_AWBURST <= twiddle_h_rsc_0_2_AWBURST;
  twiddle_h_rsc_0_2_i_AWCACHE <= twiddle_h_rsc_0_2_AWCACHE;
  twiddle_h_rsc_0_2_i_AWPROT <= twiddle_h_rsc_0_2_AWPROT;
  twiddle_h_rsc_0_2_i_AWQOS <= twiddle_h_rsc_0_2_AWQOS;
  twiddle_h_rsc_0_2_i_AWREGION <= twiddle_h_rsc_0_2_AWREGION;
  twiddle_h_rsc_0_2_i_AWUSER(0) <= twiddle_h_rsc_0_2_AWUSER;
  twiddle_h_rsc_0_2_i_WDATA <= twiddle_h_rsc_0_2_WDATA;
  twiddle_h_rsc_0_2_i_WSTRB <= twiddle_h_rsc_0_2_WSTRB;
  twiddle_h_rsc_0_2_i_WUSER(0) <= twiddle_h_rsc_0_2_WUSER;
  twiddle_h_rsc_0_2_BID <= twiddle_h_rsc_0_2_i_BID(0);
  twiddle_h_rsc_0_2_BRESP <= twiddle_h_rsc_0_2_i_BRESP;
  twiddle_h_rsc_0_2_BUSER <= twiddle_h_rsc_0_2_i_BUSER(0);
  twiddle_h_rsc_0_2_i_ARID(0) <= twiddle_h_rsc_0_2_ARID;
  twiddle_h_rsc_0_2_i_ARADDR <= twiddle_h_rsc_0_2_ARADDR;
  twiddle_h_rsc_0_2_i_ARLEN <= twiddle_h_rsc_0_2_ARLEN;
  twiddle_h_rsc_0_2_i_ARSIZE <= twiddle_h_rsc_0_2_ARSIZE;
  twiddle_h_rsc_0_2_i_ARBURST <= twiddle_h_rsc_0_2_ARBURST;
  twiddle_h_rsc_0_2_i_ARCACHE <= twiddle_h_rsc_0_2_ARCACHE;
  twiddle_h_rsc_0_2_i_ARPROT <= twiddle_h_rsc_0_2_ARPROT;
  twiddle_h_rsc_0_2_i_ARQOS <= twiddle_h_rsc_0_2_ARQOS;
  twiddle_h_rsc_0_2_i_ARREGION <= twiddle_h_rsc_0_2_ARREGION;
  twiddle_h_rsc_0_2_i_ARUSER(0) <= twiddle_h_rsc_0_2_ARUSER;
  twiddle_h_rsc_0_2_RID <= twiddle_h_rsc_0_2_i_RID(0);
  twiddle_h_rsc_0_2_RDATA <= twiddle_h_rsc_0_2_i_RDATA;
  twiddle_h_rsc_0_2_RRESP <= twiddle_h_rsc_0_2_i_RRESP;
  twiddle_h_rsc_0_2_RUSER <= twiddle_h_rsc_0_2_i_RUSER(0);
  twiddle_h_rsc_0_2_i_s_raddr_1 <= twiddle_h_rsc_0_2_i_s_raddr;
  twiddle_h_rsc_0_2_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_2_i_s_din <= twiddle_h_rsc_0_2_i_s_din_1;
  twiddle_h_rsc_0_2_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_2_i_oswt => twiddle_h_rsc_0_2_i_oswt,
      twiddle_h_rsc_0_2_i_biwt => twiddle_h_rsc_0_2_i_biwt,
      twiddle_h_rsc_0_2_i_bdwt => twiddle_h_rsc_0_2_i_bdwt,
      twiddle_h_rsc_0_2_i_bcwt => twiddle_h_rsc_0_2_i_bcwt,
      twiddle_h_rsc_0_2_i_s_re_core_sct => twiddle_h_rsc_0_2_i_s_re_core_sct,
      twiddle_h_rsc_0_2_i_s_rrdy => twiddle_h_rsc_0_2_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_2_i_oswt => twiddle_h_rsc_0_2_i_oswt,
      twiddle_h_rsc_0_2_i_wen_comp => twiddle_h_rsc_0_2_i_wen_comp,
      twiddle_h_rsc_0_2_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_s_raddr_core,
      twiddle_h_rsc_0_2_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_s_din_mxwt,
      twiddle_h_rsc_0_2_i_biwt => twiddle_h_rsc_0_2_i_biwt,
      twiddle_h_rsc_0_2_i_bdwt => twiddle_h_rsc_0_2_i_bdwt,
      twiddle_h_rsc_0_2_i_bcwt => twiddle_h_rsc_0_2_i_bcwt,
      twiddle_h_rsc_0_2_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_s_raddr,
      twiddle_h_rsc_0_2_i_s_raddr_core_sct => twiddle_h_rsc_0_2_i_s_re_core_sct,
      twiddle_h_rsc_0_2_i_s_din => peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_2_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_2_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_s_din_mxwt;
  twiddle_h_rsc_0_2_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_2_i_twiddle_h_rsc_0_2_wait_dp_inst_twiddle_h_rsc_0_2_i_s_din
      <= twiddle_h_rsc_0_2_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_1_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_1_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_1_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_1_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_1_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_1_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_1_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_1_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_1_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_1_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_1_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_1_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_1_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_1_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_1_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_1_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_1_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_1_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_1_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_1_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_1_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_1_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_1_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_1_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_1_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_1_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_1_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_1_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_1_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_1_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_1_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_1_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_1_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_1_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_1_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_1_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_1_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_1_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_1_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_1_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_1_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_1_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_1_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_1_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_1_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_1_i_AWID,
      AWADDR => twiddle_h_rsc_0_1_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_1_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_1_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_1_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_1_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_1_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_1_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_1_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_1_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_1_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_1_AWVALID,
      AWREADY => twiddle_h_rsc_0_1_AWREADY,
      WDATA => twiddle_h_rsc_0_1_i_WDATA,
      WSTRB => twiddle_h_rsc_0_1_i_WSTRB,
      WLAST => twiddle_h_rsc_0_1_WLAST,
      WUSER => twiddle_h_rsc_0_1_i_WUSER,
      WVALID => twiddle_h_rsc_0_1_WVALID,
      WREADY => twiddle_h_rsc_0_1_WREADY,
      BID => twiddle_h_rsc_0_1_i_BID,
      BRESP => twiddle_h_rsc_0_1_i_BRESP,
      BUSER => twiddle_h_rsc_0_1_i_BUSER,
      BVALID => twiddle_h_rsc_0_1_BVALID,
      BREADY => twiddle_h_rsc_0_1_BREADY,
      ARID => twiddle_h_rsc_0_1_i_ARID,
      ARADDR => twiddle_h_rsc_0_1_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_1_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_1_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_1_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_1_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_1_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_1_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_1_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_1_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_1_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_1_ARVALID,
      ARREADY => twiddle_h_rsc_0_1_ARREADY,
      RID => twiddle_h_rsc_0_1_i_RID,
      RDATA => twiddle_h_rsc_0_1_i_RDATA,
      RRESP => twiddle_h_rsc_0_1_i_RRESP,
      RLAST => twiddle_h_rsc_0_1_RLAST,
      RUSER => twiddle_h_rsc_0_1_i_RUSER,
      RVALID => twiddle_h_rsc_0_1_RVALID,
      RREADY => twiddle_h_rsc_0_1_RREADY,
      s_re => twiddle_h_rsc_0_1_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_1_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_1_i_s_waddr,
      s_din => twiddle_h_rsc_0_1_i_s_din_1,
      s_dout => twiddle_h_rsc_0_1_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_1_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_1_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_1_is_idle,
      tr_write_done => twiddle_h_rsc_0_1_tr_write_done,
      s_tdone => twiddle_h_rsc_0_1_s_tdone
    );
  twiddle_h_rsc_0_1_i_AWID(0) <= twiddle_h_rsc_0_1_AWID;
  twiddle_h_rsc_0_1_i_AWADDR <= twiddle_h_rsc_0_1_AWADDR;
  twiddle_h_rsc_0_1_i_AWLEN <= twiddle_h_rsc_0_1_AWLEN;
  twiddle_h_rsc_0_1_i_AWSIZE <= twiddle_h_rsc_0_1_AWSIZE;
  twiddle_h_rsc_0_1_i_AWBURST <= twiddle_h_rsc_0_1_AWBURST;
  twiddle_h_rsc_0_1_i_AWCACHE <= twiddle_h_rsc_0_1_AWCACHE;
  twiddle_h_rsc_0_1_i_AWPROT <= twiddle_h_rsc_0_1_AWPROT;
  twiddle_h_rsc_0_1_i_AWQOS <= twiddle_h_rsc_0_1_AWQOS;
  twiddle_h_rsc_0_1_i_AWREGION <= twiddle_h_rsc_0_1_AWREGION;
  twiddle_h_rsc_0_1_i_AWUSER(0) <= twiddle_h_rsc_0_1_AWUSER;
  twiddle_h_rsc_0_1_i_WDATA <= twiddle_h_rsc_0_1_WDATA;
  twiddle_h_rsc_0_1_i_WSTRB <= twiddle_h_rsc_0_1_WSTRB;
  twiddle_h_rsc_0_1_i_WUSER(0) <= twiddle_h_rsc_0_1_WUSER;
  twiddle_h_rsc_0_1_BID <= twiddle_h_rsc_0_1_i_BID(0);
  twiddle_h_rsc_0_1_BRESP <= twiddle_h_rsc_0_1_i_BRESP;
  twiddle_h_rsc_0_1_BUSER <= twiddle_h_rsc_0_1_i_BUSER(0);
  twiddle_h_rsc_0_1_i_ARID(0) <= twiddle_h_rsc_0_1_ARID;
  twiddle_h_rsc_0_1_i_ARADDR <= twiddle_h_rsc_0_1_ARADDR;
  twiddle_h_rsc_0_1_i_ARLEN <= twiddle_h_rsc_0_1_ARLEN;
  twiddle_h_rsc_0_1_i_ARSIZE <= twiddle_h_rsc_0_1_ARSIZE;
  twiddle_h_rsc_0_1_i_ARBURST <= twiddle_h_rsc_0_1_ARBURST;
  twiddle_h_rsc_0_1_i_ARCACHE <= twiddle_h_rsc_0_1_ARCACHE;
  twiddle_h_rsc_0_1_i_ARPROT <= twiddle_h_rsc_0_1_ARPROT;
  twiddle_h_rsc_0_1_i_ARQOS <= twiddle_h_rsc_0_1_ARQOS;
  twiddle_h_rsc_0_1_i_ARREGION <= twiddle_h_rsc_0_1_ARREGION;
  twiddle_h_rsc_0_1_i_ARUSER(0) <= twiddle_h_rsc_0_1_ARUSER;
  twiddle_h_rsc_0_1_RID <= twiddle_h_rsc_0_1_i_RID(0);
  twiddle_h_rsc_0_1_RDATA <= twiddle_h_rsc_0_1_i_RDATA;
  twiddle_h_rsc_0_1_RRESP <= twiddle_h_rsc_0_1_i_RRESP;
  twiddle_h_rsc_0_1_RUSER <= twiddle_h_rsc_0_1_i_RUSER(0);
  twiddle_h_rsc_0_1_i_s_raddr_1 <= twiddle_h_rsc_0_1_i_s_raddr;
  twiddle_h_rsc_0_1_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_1_i_s_din <= twiddle_h_rsc_0_1_i_s_din_1;
  twiddle_h_rsc_0_1_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_1_i_oswt => twiddle_h_rsc_0_1_i_oswt,
      twiddle_h_rsc_0_1_i_biwt => twiddle_h_rsc_0_1_i_biwt,
      twiddle_h_rsc_0_1_i_bdwt => twiddle_h_rsc_0_1_i_bdwt,
      twiddle_h_rsc_0_1_i_bcwt => twiddle_h_rsc_0_1_i_bcwt,
      twiddle_h_rsc_0_1_i_s_re_core_sct => twiddle_h_rsc_0_1_i_s_re_core_sct,
      twiddle_h_rsc_0_1_i_s_rrdy => twiddle_h_rsc_0_1_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_1_i_oswt => twiddle_h_rsc_0_1_i_oswt,
      twiddle_h_rsc_0_1_i_wen_comp => twiddle_h_rsc_0_1_i_wen_comp,
      twiddle_h_rsc_0_1_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_s_raddr_core,
      twiddle_h_rsc_0_1_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_s_din_mxwt,
      twiddle_h_rsc_0_1_i_biwt => twiddle_h_rsc_0_1_i_biwt,
      twiddle_h_rsc_0_1_i_bdwt => twiddle_h_rsc_0_1_i_bdwt,
      twiddle_h_rsc_0_1_i_bcwt => twiddle_h_rsc_0_1_i_bcwt,
      twiddle_h_rsc_0_1_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_s_raddr,
      twiddle_h_rsc_0_1_i_s_raddr_core_sct => twiddle_h_rsc_0_1_i_s_re_core_sct,
      twiddle_h_rsc_0_1_i_s_din => peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_1_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_1_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_s_din_mxwt;
  twiddle_h_rsc_0_1_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_1_i_twiddle_h_rsc_0_1_wait_dp_inst_twiddle_h_rsc_0_1_i_s_din
      <= twiddle_h_rsc_0_1_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_h_rsc_0_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_h_rsc_0_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_h_rsc_0_0_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_0_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_0_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_0_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_0_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_0_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_0_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_0_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_0_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_0_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_0_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_0_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_oswt : IN STD_LOGIC;
    twiddle_h_rsc_0_0_i_wen_comp : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_h_rsc_0_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_h_rsc_0_0_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_h_rsc_0_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_h_rsc_0_0_i_biwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_0_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_0_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_0_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_0_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_0_is_idle : STD_LOGIC;

  SIGNAL twiddle_h_rsc_0_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_biwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_i_bdwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_i_bcwt : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_0_i_biwt : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_bdwt : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_bcwt : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_0_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_h_rsc_0_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_h_rsc_0_0_i_AWID,
      AWADDR => twiddle_h_rsc_0_0_i_AWADDR,
      AWLEN => twiddle_h_rsc_0_0_i_AWLEN,
      AWSIZE => twiddle_h_rsc_0_0_i_AWSIZE,
      AWBURST => twiddle_h_rsc_0_0_i_AWBURST,
      AWLOCK => twiddle_h_rsc_0_0_AWLOCK,
      AWCACHE => twiddle_h_rsc_0_0_i_AWCACHE,
      AWPROT => twiddle_h_rsc_0_0_i_AWPROT,
      AWQOS => twiddle_h_rsc_0_0_i_AWQOS,
      AWREGION => twiddle_h_rsc_0_0_i_AWREGION,
      AWUSER => twiddle_h_rsc_0_0_i_AWUSER,
      AWVALID => twiddle_h_rsc_0_0_AWVALID,
      AWREADY => twiddle_h_rsc_0_0_AWREADY,
      WDATA => twiddle_h_rsc_0_0_i_WDATA,
      WSTRB => twiddle_h_rsc_0_0_i_WSTRB,
      WLAST => twiddle_h_rsc_0_0_WLAST,
      WUSER => twiddle_h_rsc_0_0_i_WUSER,
      WVALID => twiddle_h_rsc_0_0_WVALID,
      WREADY => twiddle_h_rsc_0_0_WREADY,
      BID => twiddle_h_rsc_0_0_i_BID,
      BRESP => twiddle_h_rsc_0_0_i_BRESP,
      BUSER => twiddle_h_rsc_0_0_i_BUSER,
      BVALID => twiddle_h_rsc_0_0_BVALID,
      BREADY => twiddle_h_rsc_0_0_BREADY,
      ARID => twiddle_h_rsc_0_0_i_ARID,
      ARADDR => twiddle_h_rsc_0_0_i_ARADDR,
      ARLEN => twiddle_h_rsc_0_0_i_ARLEN,
      ARSIZE => twiddle_h_rsc_0_0_i_ARSIZE,
      ARBURST => twiddle_h_rsc_0_0_i_ARBURST,
      ARLOCK => twiddle_h_rsc_0_0_ARLOCK,
      ARCACHE => twiddle_h_rsc_0_0_i_ARCACHE,
      ARPROT => twiddle_h_rsc_0_0_i_ARPROT,
      ARQOS => twiddle_h_rsc_0_0_i_ARQOS,
      ARREGION => twiddle_h_rsc_0_0_i_ARREGION,
      ARUSER => twiddle_h_rsc_0_0_i_ARUSER,
      ARVALID => twiddle_h_rsc_0_0_ARVALID,
      ARREADY => twiddle_h_rsc_0_0_ARREADY,
      RID => twiddle_h_rsc_0_0_i_RID,
      RDATA => twiddle_h_rsc_0_0_i_RDATA,
      RRESP => twiddle_h_rsc_0_0_i_RRESP,
      RLAST => twiddle_h_rsc_0_0_RLAST,
      RUSER => twiddle_h_rsc_0_0_i_RUSER,
      RVALID => twiddle_h_rsc_0_0_RVALID,
      RREADY => twiddle_h_rsc_0_0_RREADY,
      s_re => twiddle_h_rsc_0_0_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_h_rsc_0_0_i_s_raddr_1,
      s_waddr => twiddle_h_rsc_0_0_i_s_waddr,
      s_din => twiddle_h_rsc_0_0_i_s_din_1,
      s_dout => twiddle_h_rsc_0_0_i_s_dout,
      s_rrdy => twiddle_h_rsc_0_0_i_s_rrdy,
      s_wrdy => twiddle_h_rsc_0_0_i_s_wrdy,
      is_idle => twiddle_h_rsc_0_0_is_idle,
      tr_write_done => twiddle_h_rsc_0_0_tr_write_done,
      s_tdone => twiddle_h_rsc_0_0_s_tdone
    );
  twiddle_h_rsc_0_0_i_AWID(0) <= twiddle_h_rsc_0_0_AWID;
  twiddle_h_rsc_0_0_i_AWADDR <= twiddle_h_rsc_0_0_AWADDR;
  twiddle_h_rsc_0_0_i_AWLEN <= twiddle_h_rsc_0_0_AWLEN;
  twiddle_h_rsc_0_0_i_AWSIZE <= twiddle_h_rsc_0_0_AWSIZE;
  twiddle_h_rsc_0_0_i_AWBURST <= twiddle_h_rsc_0_0_AWBURST;
  twiddle_h_rsc_0_0_i_AWCACHE <= twiddle_h_rsc_0_0_AWCACHE;
  twiddle_h_rsc_0_0_i_AWPROT <= twiddle_h_rsc_0_0_AWPROT;
  twiddle_h_rsc_0_0_i_AWQOS <= twiddle_h_rsc_0_0_AWQOS;
  twiddle_h_rsc_0_0_i_AWREGION <= twiddle_h_rsc_0_0_AWREGION;
  twiddle_h_rsc_0_0_i_AWUSER(0) <= twiddle_h_rsc_0_0_AWUSER;
  twiddle_h_rsc_0_0_i_WDATA <= twiddle_h_rsc_0_0_WDATA;
  twiddle_h_rsc_0_0_i_WSTRB <= twiddle_h_rsc_0_0_WSTRB;
  twiddle_h_rsc_0_0_i_WUSER(0) <= twiddle_h_rsc_0_0_WUSER;
  twiddle_h_rsc_0_0_BID <= twiddle_h_rsc_0_0_i_BID(0);
  twiddle_h_rsc_0_0_BRESP <= twiddle_h_rsc_0_0_i_BRESP;
  twiddle_h_rsc_0_0_BUSER <= twiddle_h_rsc_0_0_i_BUSER(0);
  twiddle_h_rsc_0_0_i_ARID(0) <= twiddle_h_rsc_0_0_ARID;
  twiddle_h_rsc_0_0_i_ARADDR <= twiddle_h_rsc_0_0_ARADDR;
  twiddle_h_rsc_0_0_i_ARLEN <= twiddle_h_rsc_0_0_ARLEN;
  twiddle_h_rsc_0_0_i_ARSIZE <= twiddle_h_rsc_0_0_ARSIZE;
  twiddle_h_rsc_0_0_i_ARBURST <= twiddle_h_rsc_0_0_ARBURST;
  twiddle_h_rsc_0_0_i_ARCACHE <= twiddle_h_rsc_0_0_ARCACHE;
  twiddle_h_rsc_0_0_i_ARPROT <= twiddle_h_rsc_0_0_ARPROT;
  twiddle_h_rsc_0_0_i_ARQOS <= twiddle_h_rsc_0_0_ARQOS;
  twiddle_h_rsc_0_0_i_ARREGION <= twiddle_h_rsc_0_0_ARREGION;
  twiddle_h_rsc_0_0_i_ARUSER(0) <= twiddle_h_rsc_0_0_ARUSER;
  twiddle_h_rsc_0_0_RID <= twiddle_h_rsc_0_0_i_RID(0);
  twiddle_h_rsc_0_0_RDATA <= twiddle_h_rsc_0_0_i_RDATA;
  twiddle_h_rsc_0_0_RRESP <= twiddle_h_rsc_0_0_i_RRESP;
  twiddle_h_rsc_0_0_RUSER <= twiddle_h_rsc_0_0_i_RUSER(0);
  twiddle_h_rsc_0_0_i_s_raddr_1 <= twiddle_h_rsc_0_0_i_s_raddr;
  twiddle_h_rsc_0_0_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_h_rsc_0_0_i_s_din <= twiddle_h_rsc_0_0_i_s_din_1;
  twiddle_h_rsc_0_0_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_ctrl_inst : peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_h_rsc_0_0_i_oswt => twiddle_h_rsc_0_0_i_oswt,
      twiddle_h_rsc_0_0_i_biwt => twiddle_h_rsc_0_0_i_biwt,
      twiddle_h_rsc_0_0_i_bdwt => twiddle_h_rsc_0_0_i_bdwt,
      twiddle_h_rsc_0_0_i_bcwt => twiddle_h_rsc_0_0_i_bcwt,
      twiddle_h_rsc_0_0_i_s_re_core_sct => twiddle_h_rsc_0_0_i_s_re_core_sct,
      twiddle_h_rsc_0_0_i_s_rrdy => twiddle_h_rsc_0_0_i_s_rrdy
    );
  peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp_inst : peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_0_i_oswt => twiddle_h_rsc_0_0_i_oswt,
      twiddle_h_rsc_0_0_i_wen_comp => twiddle_h_rsc_0_0_i_wen_comp,
      twiddle_h_rsc_0_0_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_s_raddr_core,
      twiddle_h_rsc_0_0_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_s_din_mxwt,
      twiddle_h_rsc_0_0_i_biwt => twiddle_h_rsc_0_0_i_biwt,
      twiddle_h_rsc_0_0_i_bdwt => twiddle_h_rsc_0_0_i_bdwt,
      twiddle_h_rsc_0_0_i_bcwt => twiddle_h_rsc_0_0_i_bcwt,
      twiddle_h_rsc_0_0_i_s_raddr => peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_s_raddr,
      twiddle_h_rsc_0_0_i_s_raddr_core_sct => twiddle_h_rsc_0_0_i_s_re_core_sct,
      twiddle_h_rsc_0_0_i_s_din => peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_s_din
    );
  peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_s_raddr_core
      <= '0' & (twiddle_h_rsc_0_0_i_s_raddr_core(4 DOWNTO 0));
  twiddle_h_rsc_0_0_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_s_din_mxwt;
  twiddle_h_rsc_0_0_i_s_raddr <= peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_s_raddr;
  peaseNTT_core_twiddle_h_rsc_0_0_i_twiddle_h_rsc_0_0_wait_dp_inst_twiddle_h_rsc_0_0_i_s_din
      <= twiddle_h_rsc_0_0_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_15_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_15_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_15_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_15_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_15_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_15_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_15_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_15_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_15_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_15_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_15_RID : OUT STD_LOGIC;
    twiddle_rsc_0_15_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_15_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_15_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_15_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_15_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_15_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_15_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_15_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_15_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_15_ARID : IN STD_LOGIC;
    twiddle_rsc_0_15_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_15_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_15_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_15_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_15_BID : OUT STD_LOGIC;
    twiddle_rsc_0_15_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_15_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_15_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_15_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_15_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_15_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_15_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_15_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_15_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_15_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_15_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_15_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_15_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_15_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_15_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_15_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_15_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_15_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_15_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_15_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_15_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_15_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_15_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_15_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_15_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_15_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_15_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_15_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_15_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_15_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_15_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_15_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_15_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_15_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_15_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_15_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_15_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_15_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_15_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_15_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_15_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_15_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_15_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_15_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_15_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp_inst_twiddle_rsc_0_15_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp_inst_twiddle_rsc_0_15_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp_inst_twiddle_rsc_0_15_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp_inst_twiddle_rsc_0_15_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_15_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_15_i_AWID,
      AWADDR => twiddle_rsc_0_15_i_AWADDR,
      AWLEN => twiddle_rsc_0_15_i_AWLEN,
      AWSIZE => twiddle_rsc_0_15_i_AWSIZE,
      AWBURST => twiddle_rsc_0_15_i_AWBURST,
      AWLOCK => twiddle_rsc_0_15_AWLOCK,
      AWCACHE => twiddle_rsc_0_15_i_AWCACHE,
      AWPROT => twiddle_rsc_0_15_i_AWPROT,
      AWQOS => twiddle_rsc_0_15_i_AWQOS,
      AWREGION => twiddle_rsc_0_15_i_AWREGION,
      AWUSER => twiddle_rsc_0_15_i_AWUSER,
      AWVALID => twiddle_rsc_0_15_AWVALID,
      AWREADY => twiddle_rsc_0_15_AWREADY,
      WDATA => twiddle_rsc_0_15_i_WDATA,
      WSTRB => twiddle_rsc_0_15_i_WSTRB,
      WLAST => twiddle_rsc_0_15_WLAST,
      WUSER => twiddle_rsc_0_15_i_WUSER,
      WVALID => twiddle_rsc_0_15_WVALID,
      WREADY => twiddle_rsc_0_15_WREADY,
      BID => twiddle_rsc_0_15_i_BID,
      BRESP => twiddle_rsc_0_15_i_BRESP,
      BUSER => twiddle_rsc_0_15_i_BUSER,
      BVALID => twiddle_rsc_0_15_BVALID,
      BREADY => twiddle_rsc_0_15_BREADY,
      ARID => twiddle_rsc_0_15_i_ARID,
      ARADDR => twiddle_rsc_0_15_i_ARADDR,
      ARLEN => twiddle_rsc_0_15_i_ARLEN,
      ARSIZE => twiddle_rsc_0_15_i_ARSIZE,
      ARBURST => twiddle_rsc_0_15_i_ARBURST,
      ARLOCK => twiddle_rsc_0_15_ARLOCK,
      ARCACHE => twiddle_rsc_0_15_i_ARCACHE,
      ARPROT => twiddle_rsc_0_15_i_ARPROT,
      ARQOS => twiddle_rsc_0_15_i_ARQOS,
      ARREGION => twiddle_rsc_0_15_i_ARREGION,
      ARUSER => twiddle_rsc_0_15_i_ARUSER,
      ARVALID => twiddle_rsc_0_15_ARVALID,
      ARREADY => twiddle_rsc_0_15_ARREADY,
      RID => twiddle_rsc_0_15_i_RID,
      RDATA => twiddle_rsc_0_15_i_RDATA,
      RRESP => twiddle_rsc_0_15_i_RRESP,
      RLAST => twiddle_rsc_0_15_RLAST,
      RUSER => twiddle_rsc_0_15_i_RUSER,
      RVALID => twiddle_rsc_0_15_RVALID,
      RREADY => twiddle_rsc_0_15_RREADY,
      s_re => twiddle_rsc_0_15_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_15_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_15_i_s_waddr,
      s_din => twiddle_rsc_0_15_i_s_din_1,
      s_dout => twiddle_rsc_0_15_i_s_dout,
      s_rrdy => twiddle_rsc_0_15_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_15_i_s_wrdy,
      is_idle => twiddle_rsc_0_15_is_idle,
      tr_write_done => twiddle_rsc_0_15_tr_write_done,
      s_tdone => twiddle_rsc_0_15_s_tdone
    );
  twiddle_rsc_0_15_i_AWID(0) <= twiddle_rsc_0_15_AWID;
  twiddle_rsc_0_15_i_AWADDR <= twiddle_rsc_0_15_AWADDR;
  twiddle_rsc_0_15_i_AWLEN <= twiddle_rsc_0_15_AWLEN;
  twiddle_rsc_0_15_i_AWSIZE <= twiddle_rsc_0_15_AWSIZE;
  twiddle_rsc_0_15_i_AWBURST <= twiddle_rsc_0_15_AWBURST;
  twiddle_rsc_0_15_i_AWCACHE <= twiddle_rsc_0_15_AWCACHE;
  twiddle_rsc_0_15_i_AWPROT <= twiddle_rsc_0_15_AWPROT;
  twiddle_rsc_0_15_i_AWQOS <= twiddle_rsc_0_15_AWQOS;
  twiddle_rsc_0_15_i_AWREGION <= twiddle_rsc_0_15_AWREGION;
  twiddle_rsc_0_15_i_AWUSER(0) <= twiddle_rsc_0_15_AWUSER;
  twiddle_rsc_0_15_i_WDATA <= twiddle_rsc_0_15_WDATA;
  twiddle_rsc_0_15_i_WSTRB <= twiddle_rsc_0_15_WSTRB;
  twiddle_rsc_0_15_i_WUSER(0) <= twiddle_rsc_0_15_WUSER;
  twiddle_rsc_0_15_BID <= twiddle_rsc_0_15_i_BID(0);
  twiddle_rsc_0_15_BRESP <= twiddle_rsc_0_15_i_BRESP;
  twiddle_rsc_0_15_BUSER <= twiddle_rsc_0_15_i_BUSER(0);
  twiddle_rsc_0_15_i_ARID(0) <= twiddle_rsc_0_15_ARID;
  twiddle_rsc_0_15_i_ARADDR <= twiddle_rsc_0_15_ARADDR;
  twiddle_rsc_0_15_i_ARLEN <= twiddle_rsc_0_15_ARLEN;
  twiddle_rsc_0_15_i_ARSIZE <= twiddle_rsc_0_15_ARSIZE;
  twiddle_rsc_0_15_i_ARBURST <= twiddle_rsc_0_15_ARBURST;
  twiddle_rsc_0_15_i_ARCACHE <= twiddle_rsc_0_15_ARCACHE;
  twiddle_rsc_0_15_i_ARPROT <= twiddle_rsc_0_15_ARPROT;
  twiddle_rsc_0_15_i_ARQOS <= twiddle_rsc_0_15_ARQOS;
  twiddle_rsc_0_15_i_ARREGION <= twiddle_rsc_0_15_ARREGION;
  twiddle_rsc_0_15_i_ARUSER(0) <= twiddle_rsc_0_15_ARUSER;
  twiddle_rsc_0_15_RID <= twiddle_rsc_0_15_i_RID(0);
  twiddle_rsc_0_15_RDATA <= twiddle_rsc_0_15_i_RDATA;
  twiddle_rsc_0_15_RRESP <= twiddle_rsc_0_15_i_RRESP;
  twiddle_rsc_0_15_RUSER <= twiddle_rsc_0_15_i_RUSER(0);
  twiddle_rsc_0_15_i_s_raddr_1 <= twiddle_rsc_0_15_i_s_raddr;
  twiddle_rsc_0_15_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_15_i_s_din <= twiddle_rsc_0_15_i_s_din_1;
  twiddle_rsc_0_15_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_15_i_oswt => twiddle_rsc_0_15_i_oswt,
      twiddle_rsc_0_15_i_biwt => twiddle_rsc_0_15_i_biwt,
      twiddle_rsc_0_15_i_bdwt => twiddle_rsc_0_15_i_bdwt,
      twiddle_rsc_0_15_i_bcwt => twiddle_rsc_0_15_i_bcwt,
      twiddle_rsc_0_15_i_s_re_core_sct => twiddle_rsc_0_15_i_s_re_core_sct,
      twiddle_rsc_0_15_i_s_rrdy => twiddle_rsc_0_15_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_15_i_oswt => twiddle_rsc_0_15_i_oswt,
      twiddle_rsc_0_15_i_wen_comp => twiddle_rsc_0_15_i_wen_comp,
      twiddle_rsc_0_15_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp_inst_twiddle_rsc_0_15_i_s_raddr_core,
      twiddle_rsc_0_15_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp_inst_twiddle_rsc_0_15_i_s_din_mxwt,
      twiddle_rsc_0_15_i_biwt => twiddle_rsc_0_15_i_biwt,
      twiddle_rsc_0_15_i_bdwt => twiddle_rsc_0_15_i_bdwt,
      twiddle_rsc_0_15_i_bcwt => twiddle_rsc_0_15_i_bcwt,
      twiddle_rsc_0_15_i_s_raddr => peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp_inst_twiddle_rsc_0_15_i_s_raddr,
      twiddle_rsc_0_15_i_s_raddr_core_sct => twiddle_rsc_0_15_i_s_re_core_sct,
      twiddle_rsc_0_15_i_s_din => peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp_inst_twiddle_rsc_0_15_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp_inst_twiddle_rsc_0_15_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_15_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_15_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp_inst_twiddle_rsc_0_15_i_s_din_mxwt;
  twiddle_rsc_0_15_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp_inst_twiddle_rsc_0_15_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_15_i_twiddle_rsc_0_15_wait_dp_inst_twiddle_rsc_0_15_i_s_din
      <= twiddle_rsc_0_15_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_14_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_14_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_14_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_14_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_14_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_14_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_14_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_14_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_14_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_14_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_14_RID : OUT STD_LOGIC;
    twiddle_rsc_0_14_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_14_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_14_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_14_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_14_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_14_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_14_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_14_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_14_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_14_ARID : IN STD_LOGIC;
    twiddle_rsc_0_14_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_14_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_14_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_14_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_14_BID : OUT STD_LOGIC;
    twiddle_rsc_0_14_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_14_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_14_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_14_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_14_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_14_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_14_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_14_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_14_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_14_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_14_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_14_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_14_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_14_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_14_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_14_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_14_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_14_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_14_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_14_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_14_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_14_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_14_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_14_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_14_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_14_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_14_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_14_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_14_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_14_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_14_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_14_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_14_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_14_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_14_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_14_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_14_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_14_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_14_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_14_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_14_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_14_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_14_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_14_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_14_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp_inst_twiddle_rsc_0_14_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp_inst_twiddle_rsc_0_14_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp_inst_twiddle_rsc_0_14_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp_inst_twiddle_rsc_0_14_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_14_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_14_i_AWID,
      AWADDR => twiddle_rsc_0_14_i_AWADDR,
      AWLEN => twiddle_rsc_0_14_i_AWLEN,
      AWSIZE => twiddle_rsc_0_14_i_AWSIZE,
      AWBURST => twiddle_rsc_0_14_i_AWBURST,
      AWLOCK => twiddle_rsc_0_14_AWLOCK,
      AWCACHE => twiddle_rsc_0_14_i_AWCACHE,
      AWPROT => twiddle_rsc_0_14_i_AWPROT,
      AWQOS => twiddle_rsc_0_14_i_AWQOS,
      AWREGION => twiddle_rsc_0_14_i_AWREGION,
      AWUSER => twiddle_rsc_0_14_i_AWUSER,
      AWVALID => twiddle_rsc_0_14_AWVALID,
      AWREADY => twiddle_rsc_0_14_AWREADY,
      WDATA => twiddle_rsc_0_14_i_WDATA,
      WSTRB => twiddle_rsc_0_14_i_WSTRB,
      WLAST => twiddle_rsc_0_14_WLAST,
      WUSER => twiddle_rsc_0_14_i_WUSER,
      WVALID => twiddle_rsc_0_14_WVALID,
      WREADY => twiddle_rsc_0_14_WREADY,
      BID => twiddle_rsc_0_14_i_BID,
      BRESP => twiddle_rsc_0_14_i_BRESP,
      BUSER => twiddle_rsc_0_14_i_BUSER,
      BVALID => twiddle_rsc_0_14_BVALID,
      BREADY => twiddle_rsc_0_14_BREADY,
      ARID => twiddle_rsc_0_14_i_ARID,
      ARADDR => twiddle_rsc_0_14_i_ARADDR,
      ARLEN => twiddle_rsc_0_14_i_ARLEN,
      ARSIZE => twiddle_rsc_0_14_i_ARSIZE,
      ARBURST => twiddle_rsc_0_14_i_ARBURST,
      ARLOCK => twiddle_rsc_0_14_ARLOCK,
      ARCACHE => twiddle_rsc_0_14_i_ARCACHE,
      ARPROT => twiddle_rsc_0_14_i_ARPROT,
      ARQOS => twiddle_rsc_0_14_i_ARQOS,
      ARREGION => twiddle_rsc_0_14_i_ARREGION,
      ARUSER => twiddle_rsc_0_14_i_ARUSER,
      ARVALID => twiddle_rsc_0_14_ARVALID,
      ARREADY => twiddle_rsc_0_14_ARREADY,
      RID => twiddle_rsc_0_14_i_RID,
      RDATA => twiddle_rsc_0_14_i_RDATA,
      RRESP => twiddle_rsc_0_14_i_RRESP,
      RLAST => twiddle_rsc_0_14_RLAST,
      RUSER => twiddle_rsc_0_14_i_RUSER,
      RVALID => twiddle_rsc_0_14_RVALID,
      RREADY => twiddle_rsc_0_14_RREADY,
      s_re => twiddle_rsc_0_14_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_14_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_14_i_s_waddr,
      s_din => twiddle_rsc_0_14_i_s_din_1,
      s_dout => twiddle_rsc_0_14_i_s_dout,
      s_rrdy => twiddle_rsc_0_14_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_14_i_s_wrdy,
      is_idle => twiddle_rsc_0_14_is_idle,
      tr_write_done => twiddle_rsc_0_14_tr_write_done,
      s_tdone => twiddle_rsc_0_14_s_tdone
    );
  twiddle_rsc_0_14_i_AWID(0) <= twiddle_rsc_0_14_AWID;
  twiddle_rsc_0_14_i_AWADDR <= twiddle_rsc_0_14_AWADDR;
  twiddle_rsc_0_14_i_AWLEN <= twiddle_rsc_0_14_AWLEN;
  twiddle_rsc_0_14_i_AWSIZE <= twiddle_rsc_0_14_AWSIZE;
  twiddle_rsc_0_14_i_AWBURST <= twiddle_rsc_0_14_AWBURST;
  twiddle_rsc_0_14_i_AWCACHE <= twiddle_rsc_0_14_AWCACHE;
  twiddle_rsc_0_14_i_AWPROT <= twiddle_rsc_0_14_AWPROT;
  twiddle_rsc_0_14_i_AWQOS <= twiddle_rsc_0_14_AWQOS;
  twiddle_rsc_0_14_i_AWREGION <= twiddle_rsc_0_14_AWREGION;
  twiddle_rsc_0_14_i_AWUSER(0) <= twiddle_rsc_0_14_AWUSER;
  twiddle_rsc_0_14_i_WDATA <= twiddle_rsc_0_14_WDATA;
  twiddle_rsc_0_14_i_WSTRB <= twiddle_rsc_0_14_WSTRB;
  twiddle_rsc_0_14_i_WUSER(0) <= twiddle_rsc_0_14_WUSER;
  twiddle_rsc_0_14_BID <= twiddle_rsc_0_14_i_BID(0);
  twiddle_rsc_0_14_BRESP <= twiddle_rsc_0_14_i_BRESP;
  twiddle_rsc_0_14_BUSER <= twiddle_rsc_0_14_i_BUSER(0);
  twiddle_rsc_0_14_i_ARID(0) <= twiddle_rsc_0_14_ARID;
  twiddle_rsc_0_14_i_ARADDR <= twiddle_rsc_0_14_ARADDR;
  twiddle_rsc_0_14_i_ARLEN <= twiddle_rsc_0_14_ARLEN;
  twiddle_rsc_0_14_i_ARSIZE <= twiddle_rsc_0_14_ARSIZE;
  twiddle_rsc_0_14_i_ARBURST <= twiddle_rsc_0_14_ARBURST;
  twiddle_rsc_0_14_i_ARCACHE <= twiddle_rsc_0_14_ARCACHE;
  twiddle_rsc_0_14_i_ARPROT <= twiddle_rsc_0_14_ARPROT;
  twiddle_rsc_0_14_i_ARQOS <= twiddle_rsc_0_14_ARQOS;
  twiddle_rsc_0_14_i_ARREGION <= twiddle_rsc_0_14_ARREGION;
  twiddle_rsc_0_14_i_ARUSER(0) <= twiddle_rsc_0_14_ARUSER;
  twiddle_rsc_0_14_RID <= twiddle_rsc_0_14_i_RID(0);
  twiddle_rsc_0_14_RDATA <= twiddle_rsc_0_14_i_RDATA;
  twiddle_rsc_0_14_RRESP <= twiddle_rsc_0_14_i_RRESP;
  twiddle_rsc_0_14_RUSER <= twiddle_rsc_0_14_i_RUSER(0);
  twiddle_rsc_0_14_i_s_raddr_1 <= twiddle_rsc_0_14_i_s_raddr;
  twiddle_rsc_0_14_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_14_i_s_din <= twiddle_rsc_0_14_i_s_din_1;
  twiddle_rsc_0_14_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_14_i_oswt => twiddle_rsc_0_14_i_oswt,
      twiddle_rsc_0_14_i_biwt => twiddle_rsc_0_14_i_biwt,
      twiddle_rsc_0_14_i_bdwt => twiddle_rsc_0_14_i_bdwt,
      twiddle_rsc_0_14_i_bcwt => twiddle_rsc_0_14_i_bcwt,
      twiddle_rsc_0_14_i_s_re_core_sct => twiddle_rsc_0_14_i_s_re_core_sct,
      twiddle_rsc_0_14_i_s_rrdy => twiddle_rsc_0_14_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_14_i_oswt => twiddle_rsc_0_14_i_oswt,
      twiddle_rsc_0_14_i_wen_comp => twiddle_rsc_0_14_i_wen_comp,
      twiddle_rsc_0_14_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp_inst_twiddle_rsc_0_14_i_s_raddr_core,
      twiddle_rsc_0_14_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp_inst_twiddle_rsc_0_14_i_s_din_mxwt,
      twiddle_rsc_0_14_i_biwt => twiddle_rsc_0_14_i_biwt,
      twiddle_rsc_0_14_i_bdwt => twiddle_rsc_0_14_i_bdwt,
      twiddle_rsc_0_14_i_bcwt => twiddle_rsc_0_14_i_bcwt,
      twiddle_rsc_0_14_i_s_raddr => peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp_inst_twiddle_rsc_0_14_i_s_raddr,
      twiddle_rsc_0_14_i_s_raddr_core_sct => twiddle_rsc_0_14_i_s_re_core_sct,
      twiddle_rsc_0_14_i_s_din => peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp_inst_twiddle_rsc_0_14_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp_inst_twiddle_rsc_0_14_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_14_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_14_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp_inst_twiddle_rsc_0_14_i_s_din_mxwt;
  twiddle_rsc_0_14_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp_inst_twiddle_rsc_0_14_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_14_i_twiddle_rsc_0_14_wait_dp_inst_twiddle_rsc_0_14_i_s_din
      <= twiddle_rsc_0_14_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_13_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_13_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_13_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_13_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_13_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_13_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_13_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_13_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_13_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_13_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_13_RID : OUT STD_LOGIC;
    twiddle_rsc_0_13_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_13_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_13_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_13_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_13_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_13_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_13_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_13_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_13_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_13_ARID : IN STD_LOGIC;
    twiddle_rsc_0_13_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_13_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_13_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_13_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_13_BID : OUT STD_LOGIC;
    twiddle_rsc_0_13_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_13_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_13_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_13_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_13_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_13_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_13_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_13_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_13_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_13_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_13_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_13_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_13_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_13_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_13_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_13_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_13_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_13_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_13_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_13_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_13_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_13_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_13_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_13_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_13_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_13_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_13_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_13_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_13_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_13_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_13_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_13_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_13_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_13_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_13_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_13_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_13_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_13_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_13_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_13_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_13_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_13_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_13_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_13_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_13_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp_inst_twiddle_rsc_0_13_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp_inst_twiddle_rsc_0_13_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp_inst_twiddle_rsc_0_13_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp_inst_twiddle_rsc_0_13_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_13_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_13_i_AWID,
      AWADDR => twiddle_rsc_0_13_i_AWADDR,
      AWLEN => twiddle_rsc_0_13_i_AWLEN,
      AWSIZE => twiddle_rsc_0_13_i_AWSIZE,
      AWBURST => twiddle_rsc_0_13_i_AWBURST,
      AWLOCK => twiddle_rsc_0_13_AWLOCK,
      AWCACHE => twiddle_rsc_0_13_i_AWCACHE,
      AWPROT => twiddle_rsc_0_13_i_AWPROT,
      AWQOS => twiddle_rsc_0_13_i_AWQOS,
      AWREGION => twiddle_rsc_0_13_i_AWREGION,
      AWUSER => twiddle_rsc_0_13_i_AWUSER,
      AWVALID => twiddle_rsc_0_13_AWVALID,
      AWREADY => twiddle_rsc_0_13_AWREADY,
      WDATA => twiddle_rsc_0_13_i_WDATA,
      WSTRB => twiddle_rsc_0_13_i_WSTRB,
      WLAST => twiddle_rsc_0_13_WLAST,
      WUSER => twiddle_rsc_0_13_i_WUSER,
      WVALID => twiddle_rsc_0_13_WVALID,
      WREADY => twiddle_rsc_0_13_WREADY,
      BID => twiddle_rsc_0_13_i_BID,
      BRESP => twiddle_rsc_0_13_i_BRESP,
      BUSER => twiddle_rsc_0_13_i_BUSER,
      BVALID => twiddle_rsc_0_13_BVALID,
      BREADY => twiddle_rsc_0_13_BREADY,
      ARID => twiddle_rsc_0_13_i_ARID,
      ARADDR => twiddle_rsc_0_13_i_ARADDR,
      ARLEN => twiddle_rsc_0_13_i_ARLEN,
      ARSIZE => twiddle_rsc_0_13_i_ARSIZE,
      ARBURST => twiddle_rsc_0_13_i_ARBURST,
      ARLOCK => twiddle_rsc_0_13_ARLOCK,
      ARCACHE => twiddle_rsc_0_13_i_ARCACHE,
      ARPROT => twiddle_rsc_0_13_i_ARPROT,
      ARQOS => twiddle_rsc_0_13_i_ARQOS,
      ARREGION => twiddle_rsc_0_13_i_ARREGION,
      ARUSER => twiddle_rsc_0_13_i_ARUSER,
      ARVALID => twiddle_rsc_0_13_ARVALID,
      ARREADY => twiddle_rsc_0_13_ARREADY,
      RID => twiddle_rsc_0_13_i_RID,
      RDATA => twiddle_rsc_0_13_i_RDATA,
      RRESP => twiddle_rsc_0_13_i_RRESP,
      RLAST => twiddle_rsc_0_13_RLAST,
      RUSER => twiddle_rsc_0_13_i_RUSER,
      RVALID => twiddle_rsc_0_13_RVALID,
      RREADY => twiddle_rsc_0_13_RREADY,
      s_re => twiddle_rsc_0_13_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_13_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_13_i_s_waddr,
      s_din => twiddle_rsc_0_13_i_s_din_1,
      s_dout => twiddle_rsc_0_13_i_s_dout,
      s_rrdy => twiddle_rsc_0_13_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_13_i_s_wrdy,
      is_idle => twiddle_rsc_0_13_is_idle,
      tr_write_done => twiddle_rsc_0_13_tr_write_done,
      s_tdone => twiddle_rsc_0_13_s_tdone
    );
  twiddle_rsc_0_13_i_AWID(0) <= twiddle_rsc_0_13_AWID;
  twiddle_rsc_0_13_i_AWADDR <= twiddle_rsc_0_13_AWADDR;
  twiddle_rsc_0_13_i_AWLEN <= twiddle_rsc_0_13_AWLEN;
  twiddle_rsc_0_13_i_AWSIZE <= twiddle_rsc_0_13_AWSIZE;
  twiddle_rsc_0_13_i_AWBURST <= twiddle_rsc_0_13_AWBURST;
  twiddle_rsc_0_13_i_AWCACHE <= twiddle_rsc_0_13_AWCACHE;
  twiddle_rsc_0_13_i_AWPROT <= twiddle_rsc_0_13_AWPROT;
  twiddle_rsc_0_13_i_AWQOS <= twiddle_rsc_0_13_AWQOS;
  twiddle_rsc_0_13_i_AWREGION <= twiddle_rsc_0_13_AWREGION;
  twiddle_rsc_0_13_i_AWUSER(0) <= twiddle_rsc_0_13_AWUSER;
  twiddle_rsc_0_13_i_WDATA <= twiddle_rsc_0_13_WDATA;
  twiddle_rsc_0_13_i_WSTRB <= twiddle_rsc_0_13_WSTRB;
  twiddle_rsc_0_13_i_WUSER(0) <= twiddle_rsc_0_13_WUSER;
  twiddle_rsc_0_13_BID <= twiddle_rsc_0_13_i_BID(0);
  twiddle_rsc_0_13_BRESP <= twiddle_rsc_0_13_i_BRESP;
  twiddle_rsc_0_13_BUSER <= twiddle_rsc_0_13_i_BUSER(0);
  twiddle_rsc_0_13_i_ARID(0) <= twiddle_rsc_0_13_ARID;
  twiddle_rsc_0_13_i_ARADDR <= twiddle_rsc_0_13_ARADDR;
  twiddle_rsc_0_13_i_ARLEN <= twiddle_rsc_0_13_ARLEN;
  twiddle_rsc_0_13_i_ARSIZE <= twiddle_rsc_0_13_ARSIZE;
  twiddle_rsc_0_13_i_ARBURST <= twiddle_rsc_0_13_ARBURST;
  twiddle_rsc_0_13_i_ARCACHE <= twiddle_rsc_0_13_ARCACHE;
  twiddle_rsc_0_13_i_ARPROT <= twiddle_rsc_0_13_ARPROT;
  twiddle_rsc_0_13_i_ARQOS <= twiddle_rsc_0_13_ARQOS;
  twiddle_rsc_0_13_i_ARREGION <= twiddle_rsc_0_13_ARREGION;
  twiddle_rsc_0_13_i_ARUSER(0) <= twiddle_rsc_0_13_ARUSER;
  twiddle_rsc_0_13_RID <= twiddle_rsc_0_13_i_RID(0);
  twiddle_rsc_0_13_RDATA <= twiddle_rsc_0_13_i_RDATA;
  twiddle_rsc_0_13_RRESP <= twiddle_rsc_0_13_i_RRESP;
  twiddle_rsc_0_13_RUSER <= twiddle_rsc_0_13_i_RUSER(0);
  twiddle_rsc_0_13_i_s_raddr_1 <= twiddle_rsc_0_13_i_s_raddr;
  twiddle_rsc_0_13_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_13_i_s_din <= twiddle_rsc_0_13_i_s_din_1;
  twiddle_rsc_0_13_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_13_i_oswt => twiddle_rsc_0_13_i_oswt,
      twiddle_rsc_0_13_i_biwt => twiddle_rsc_0_13_i_biwt,
      twiddle_rsc_0_13_i_bdwt => twiddle_rsc_0_13_i_bdwt,
      twiddle_rsc_0_13_i_bcwt => twiddle_rsc_0_13_i_bcwt,
      twiddle_rsc_0_13_i_s_re_core_sct => twiddle_rsc_0_13_i_s_re_core_sct,
      twiddle_rsc_0_13_i_s_rrdy => twiddle_rsc_0_13_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_13_i_oswt => twiddle_rsc_0_13_i_oswt,
      twiddle_rsc_0_13_i_wen_comp => twiddle_rsc_0_13_i_wen_comp,
      twiddle_rsc_0_13_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp_inst_twiddle_rsc_0_13_i_s_raddr_core,
      twiddle_rsc_0_13_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp_inst_twiddle_rsc_0_13_i_s_din_mxwt,
      twiddle_rsc_0_13_i_biwt => twiddle_rsc_0_13_i_biwt,
      twiddle_rsc_0_13_i_bdwt => twiddle_rsc_0_13_i_bdwt,
      twiddle_rsc_0_13_i_bcwt => twiddle_rsc_0_13_i_bcwt,
      twiddle_rsc_0_13_i_s_raddr => peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp_inst_twiddle_rsc_0_13_i_s_raddr,
      twiddle_rsc_0_13_i_s_raddr_core_sct => twiddle_rsc_0_13_i_s_re_core_sct,
      twiddle_rsc_0_13_i_s_din => peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp_inst_twiddle_rsc_0_13_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp_inst_twiddle_rsc_0_13_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_13_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_13_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp_inst_twiddle_rsc_0_13_i_s_din_mxwt;
  twiddle_rsc_0_13_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp_inst_twiddle_rsc_0_13_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_13_i_twiddle_rsc_0_13_wait_dp_inst_twiddle_rsc_0_13_i_s_din
      <= twiddle_rsc_0_13_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_12_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_12_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_12_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_12_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_12_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_12_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_12_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_12_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_12_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_12_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_12_RID : OUT STD_LOGIC;
    twiddle_rsc_0_12_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_12_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_12_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_12_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_12_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_12_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_12_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_12_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_12_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_12_ARID : IN STD_LOGIC;
    twiddle_rsc_0_12_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_12_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_12_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_12_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_12_BID : OUT STD_LOGIC;
    twiddle_rsc_0_12_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_12_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_12_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_12_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_12_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_12_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_12_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_12_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_12_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_12_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_12_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_12_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_12_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_12_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_12_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_12_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_12_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_12_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_12_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_12_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_12_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_12_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_12_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_12_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_12_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_12_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_12_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_12_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_12_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_12_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_12_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_12_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_12_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_12_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_12_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_12_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_12_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_12_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_12_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_12_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_12_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_12_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_12_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_12_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_12_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp_inst_twiddle_rsc_0_12_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp_inst_twiddle_rsc_0_12_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp_inst_twiddle_rsc_0_12_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp_inst_twiddle_rsc_0_12_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_12_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_12_i_AWID,
      AWADDR => twiddle_rsc_0_12_i_AWADDR,
      AWLEN => twiddle_rsc_0_12_i_AWLEN,
      AWSIZE => twiddle_rsc_0_12_i_AWSIZE,
      AWBURST => twiddle_rsc_0_12_i_AWBURST,
      AWLOCK => twiddle_rsc_0_12_AWLOCK,
      AWCACHE => twiddle_rsc_0_12_i_AWCACHE,
      AWPROT => twiddle_rsc_0_12_i_AWPROT,
      AWQOS => twiddle_rsc_0_12_i_AWQOS,
      AWREGION => twiddle_rsc_0_12_i_AWREGION,
      AWUSER => twiddle_rsc_0_12_i_AWUSER,
      AWVALID => twiddle_rsc_0_12_AWVALID,
      AWREADY => twiddle_rsc_0_12_AWREADY,
      WDATA => twiddle_rsc_0_12_i_WDATA,
      WSTRB => twiddle_rsc_0_12_i_WSTRB,
      WLAST => twiddle_rsc_0_12_WLAST,
      WUSER => twiddle_rsc_0_12_i_WUSER,
      WVALID => twiddle_rsc_0_12_WVALID,
      WREADY => twiddle_rsc_0_12_WREADY,
      BID => twiddle_rsc_0_12_i_BID,
      BRESP => twiddle_rsc_0_12_i_BRESP,
      BUSER => twiddle_rsc_0_12_i_BUSER,
      BVALID => twiddle_rsc_0_12_BVALID,
      BREADY => twiddle_rsc_0_12_BREADY,
      ARID => twiddle_rsc_0_12_i_ARID,
      ARADDR => twiddle_rsc_0_12_i_ARADDR,
      ARLEN => twiddle_rsc_0_12_i_ARLEN,
      ARSIZE => twiddle_rsc_0_12_i_ARSIZE,
      ARBURST => twiddle_rsc_0_12_i_ARBURST,
      ARLOCK => twiddle_rsc_0_12_ARLOCK,
      ARCACHE => twiddle_rsc_0_12_i_ARCACHE,
      ARPROT => twiddle_rsc_0_12_i_ARPROT,
      ARQOS => twiddle_rsc_0_12_i_ARQOS,
      ARREGION => twiddle_rsc_0_12_i_ARREGION,
      ARUSER => twiddle_rsc_0_12_i_ARUSER,
      ARVALID => twiddle_rsc_0_12_ARVALID,
      ARREADY => twiddle_rsc_0_12_ARREADY,
      RID => twiddle_rsc_0_12_i_RID,
      RDATA => twiddle_rsc_0_12_i_RDATA,
      RRESP => twiddle_rsc_0_12_i_RRESP,
      RLAST => twiddle_rsc_0_12_RLAST,
      RUSER => twiddle_rsc_0_12_i_RUSER,
      RVALID => twiddle_rsc_0_12_RVALID,
      RREADY => twiddle_rsc_0_12_RREADY,
      s_re => twiddle_rsc_0_12_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_12_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_12_i_s_waddr,
      s_din => twiddle_rsc_0_12_i_s_din_1,
      s_dout => twiddle_rsc_0_12_i_s_dout,
      s_rrdy => twiddle_rsc_0_12_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_12_i_s_wrdy,
      is_idle => twiddle_rsc_0_12_is_idle,
      tr_write_done => twiddle_rsc_0_12_tr_write_done,
      s_tdone => twiddle_rsc_0_12_s_tdone
    );
  twiddle_rsc_0_12_i_AWID(0) <= twiddle_rsc_0_12_AWID;
  twiddle_rsc_0_12_i_AWADDR <= twiddle_rsc_0_12_AWADDR;
  twiddle_rsc_0_12_i_AWLEN <= twiddle_rsc_0_12_AWLEN;
  twiddle_rsc_0_12_i_AWSIZE <= twiddle_rsc_0_12_AWSIZE;
  twiddle_rsc_0_12_i_AWBURST <= twiddle_rsc_0_12_AWBURST;
  twiddle_rsc_0_12_i_AWCACHE <= twiddle_rsc_0_12_AWCACHE;
  twiddle_rsc_0_12_i_AWPROT <= twiddle_rsc_0_12_AWPROT;
  twiddle_rsc_0_12_i_AWQOS <= twiddle_rsc_0_12_AWQOS;
  twiddle_rsc_0_12_i_AWREGION <= twiddle_rsc_0_12_AWREGION;
  twiddle_rsc_0_12_i_AWUSER(0) <= twiddle_rsc_0_12_AWUSER;
  twiddle_rsc_0_12_i_WDATA <= twiddle_rsc_0_12_WDATA;
  twiddle_rsc_0_12_i_WSTRB <= twiddle_rsc_0_12_WSTRB;
  twiddle_rsc_0_12_i_WUSER(0) <= twiddle_rsc_0_12_WUSER;
  twiddle_rsc_0_12_BID <= twiddle_rsc_0_12_i_BID(0);
  twiddle_rsc_0_12_BRESP <= twiddle_rsc_0_12_i_BRESP;
  twiddle_rsc_0_12_BUSER <= twiddle_rsc_0_12_i_BUSER(0);
  twiddle_rsc_0_12_i_ARID(0) <= twiddle_rsc_0_12_ARID;
  twiddle_rsc_0_12_i_ARADDR <= twiddle_rsc_0_12_ARADDR;
  twiddle_rsc_0_12_i_ARLEN <= twiddle_rsc_0_12_ARLEN;
  twiddle_rsc_0_12_i_ARSIZE <= twiddle_rsc_0_12_ARSIZE;
  twiddle_rsc_0_12_i_ARBURST <= twiddle_rsc_0_12_ARBURST;
  twiddle_rsc_0_12_i_ARCACHE <= twiddle_rsc_0_12_ARCACHE;
  twiddle_rsc_0_12_i_ARPROT <= twiddle_rsc_0_12_ARPROT;
  twiddle_rsc_0_12_i_ARQOS <= twiddle_rsc_0_12_ARQOS;
  twiddle_rsc_0_12_i_ARREGION <= twiddle_rsc_0_12_ARREGION;
  twiddle_rsc_0_12_i_ARUSER(0) <= twiddle_rsc_0_12_ARUSER;
  twiddle_rsc_0_12_RID <= twiddle_rsc_0_12_i_RID(0);
  twiddle_rsc_0_12_RDATA <= twiddle_rsc_0_12_i_RDATA;
  twiddle_rsc_0_12_RRESP <= twiddle_rsc_0_12_i_RRESP;
  twiddle_rsc_0_12_RUSER <= twiddle_rsc_0_12_i_RUSER(0);
  twiddle_rsc_0_12_i_s_raddr_1 <= twiddle_rsc_0_12_i_s_raddr;
  twiddle_rsc_0_12_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_12_i_s_din <= twiddle_rsc_0_12_i_s_din_1;
  twiddle_rsc_0_12_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_12_i_oswt => twiddle_rsc_0_12_i_oswt,
      twiddle_rsc_0_12_i_biwt => twiddle_rsc_0_12_i_biwt,
      twiddle_rsc_0_12_i_bdwt => twiddle_rsc_0_12_i_bdwt,
      twiddle_rsc_0_12_i_bcwt => twiddle_rsc_0_12_i_bcwt,
      twiddle_rsc_0_12_i_s_re_core_sct => twiddle_rsc_0_12_i_s_re_core_sct,
      twiddle_rsc_0_12_i_s_rrdy => twiddle_rsc_0_12_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_12_i_oswt => twiddle_rsc_0_12_i_oswt,
      twiddle_rsc_0_12_i_wen_comp => twiddle_rsc_0_12_i_wen_comp,
      twiddle_rsc_0_12_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp_inst_twiddle_rsc_0_12_i_s_raddr_core,
      twiddle_rsc_0_12_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp_inst_twiddle_rsc_0_12_i_s_din_mxwt,
      twiddle_rsc_0_12_i_biwt => twiddle_rsc_0_12_i_biwt,
      twiddle_rsc_0_12_i_bdwt => twiddle_rsc_0_12_i_bdwt,
      twiddle_rsc_0_12_i_bcwt => twiddle_rsc_0_12_i_bcwt,
      twiddle_rsc_0_12_i_s_raddr => peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp_inst_twiddle_rsc_0_12_i_s_raddr,
      twiddle_rsc_0_12_i_s_raddr_core_sct => twiddle_rsc_0_12_i_s_re_core_sct,
      twiddle_rsc_0_12_i_s_din => peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp_inst_twiddle_rsc_0_12_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp_inst_twiddle_rsc_0_12_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_12_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_12_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp_inst_twiddle_rsc_0_12_i_s_din_mxwt;
  twiddle_rsc_0_12_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp_inst_twiddle_rsc_0_12_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_12_i_twiddle_rsc_0_12_wait_dp_inst_twiddle_rsc_0_12_i_s_din
      <= twiddle_rsc_0_12_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_11_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_11_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_11_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_11_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_11_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_11_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_11_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_11_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_11_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_11_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_11_RID : OUT STD_LOGIC;
    twiddle_rsc_0_11_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_11_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_11_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_11_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_11_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_11_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_11_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_11_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_11_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_11_ARID : IN STD_LOGIC;
    twiddle_rsc_0_11_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_11_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_11_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_11_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_11_BID : OUT STD_LOGIC;
    twiddle_rsc_0_11_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_11_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_11_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_11_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_11_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_11_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_11_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_11_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_11_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_11_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_11_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_11_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_11_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_11_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_11_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_11_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_11_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_11_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_11_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_11_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_11_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_11_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_11_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_11_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_11_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_11_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_11_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_11_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_11_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_11_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_11_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_11_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_11_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_11_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_11_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_11_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_11_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_11_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_11_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_11_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_11_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_11_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_11_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_11_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_11_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp_inst_twiddle_rsc_0_11_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp_inst_twiddle_rsc_0_11_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp_inst_twiddle_rsc_0_11_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp_inst_twiddle_rsc_0_11_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_11_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_11_i_AWID,
      AWADDR => twiddle_rsc_0_11_i_AWADDR,
      AWLEN => twiddle_rsc_0_11_i_AWLEN,
      AWSIZE => twiddle_rsc_0_11_i_AWSIZE,
      AWBURST => twiddle_rsc_0_11_i_AWBURST,
      AWLOCK => twiddle_rsc_0_11_AWLOCK,
      AWCACHE => twiddle_rsc_0_11_i_AWCACHE,
      AWPROT => twiddle_rsc_0_11_i_AWPROT,
      AWQOS => twiddle_rsc_0_11_i_AWQOS,
      AWREGION => twiddle_rsc_0_11_i_AWREGION,
      AWUSER => twiddle_rsc_0_11_i_AWUSER,
      AWVALID => twiddle_rsc_0_11_AWVALID,
      AWREADY => twiddle_rsc_0_11_AWREADY,
      WDATA => twiddle_rsc_0_11_i_WDATA,
      WSTRB => twiddle_rsc_0_11_i_WSTRB,
      WLAST => twiddle_rsc_0_11_WLAST,
      WUSER => twiddle_rsc_0_11_i_WUSER,
      WVALID => twiddle_rsc_0_11_WVALID,
      WREADY => twiddle_rsc_0_11_WREADY,
      BID => twiddle_rsc_0_11_i_BID,
      BRESP => twiddle_rsc_0_11_i_BRESP,
      BUSER => twiddle_rsc_0_11_i_BUSER,
      BVALID => twiddle_rsc_0_11_BVALID,
      BREADY => twiddle_rsc_0_11_BREADY,
      ARID => twiddle_rsc_0_11_i_ARID,
      ARADDR => twiddle_rsc_0_11_i_ARADDR,
      ARLEN => twiddle_rsc_0_11_i_ARLEN,
      ARSIZE => twiddle_rsc_0_11_i_ARSIZE,
      ARBURST => twiddle_rsc_0_11_i_ARBURST,
      ARLOCK => twiddle_rsc_0_11_ARLOCK,
      ARCACHE => twiddle_rsc_0_11_i_ARCACHE,
      ARPROT => twiddle_rsc_0_11_i_ARPROT,
      ARQOS => twiddle_rsc_0_11_i_ARQOS,
      ARREGION => twiddle_rsc_0_11_i_ARREGION,
      ARUSER => twiddle_rsc_0_11_i_ARUSER,
      ARVALID => twiddle_rsc_0_11_ARVALID,
      ARREADY => twiddle_rsc_0_11_ARREADY,
      RID => twiddle_rsc_0_11_i_RID,
      RDATA => twiddle_rsc_0_11_i_RDATA,
      RRESP => twiddle_rsc_0_11_i_RRESP,
      RLAST => twiddle_rsc_0_11_RLAST,
      RUSER => twiddle_rsc_0_11_i_RUSER,
      RVALID => twiddle_rsc_0_11_RVALID,
      RREADY => twiddle_rsc_0_11_RREADY,
      s_re => twiddle_rsc_0_11_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_11_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_11_i_s_waddr,
      s_din => twiddle_rsc_0_11_i_s_din_1,
      s_dout => twiddle_rsc_0_11_i_s_dout,
      s_rrdy => twiddle_rsc_0_11_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_11_i_s_wrdy,
      is_idle => twiddle_rsc_0_11_is_idle,
      tr_write_done => twiddle_rsc_0_11_tr_write_done,
      s_tdone => twiddle_rsc_0_11_s_tdone
    );
  twiddle_rsc_0_11_i_AWID(0) <= twiddle_rsc_0_11_AWID;
  twiddle_rsc_0_11_i_AWADDR <= twiddle_rsc_0_11_AWADDR;
  twiddle_rsc_0_11_i_AWLEN <= twiddle_rsc_0_11_AWLEN;
  twiddle_rsc_0_11_i_AWSIZE <= twiddle_rsc_0_11_AWSIZE;
  twiddle_rsc_0_11_i_AWBURST <= twiddle_rsc_0_11_AWBURST;
  twiddle_rsc_0_11_i_AWCACHE <= twiddle_rsc_0_11_AWCACHE;
  twiddle_rsc_0_11_i_AWPROT <= twiddle_rsc_0_11_AWPROT;
  twiddle_rsc_0_11_i_AWQOS <= twiddle_rsc_0_11_AWQOS;
  twiddle_rsc_0_11_i_AWREGION <= twiddle_rsc_0_11_AWREGION;
  twiddle_rsc_0_11_i_AWUSER(0) <= twiddle_rsc_0_11_AWUSER;
  twiddle_rsc_0_11_i_WDATA <= twiddle_rsc_0_11_WDATA;
  twiddle_rsc_0_11_i_WSTRB <= twiddle_rsc_0_11_WSTRB;
  twiddle_rsc_0_11_i_WUSER(0) <= twiddle_rsc_0_11_WUSER;
  twiddle_rsc_0_11_BID <= twiddle_rsc_0_11_i_BID(0);
  twiddle_rsc_0_11_BRESP <= twiddle_rsc_0_11_i_BRESP;
  twiddle_rsc_0_11_BUSER <= twiddle_rsc_0_11_i_BUSER(0);
  twiddle_rsc_0_11_i_ARID(0) <= twiddle_rsc_0_11_ARID;
  twiddle_rsc_0_11_i_ARADDR <= twiddle_rsc_0_11_ARADDR;
  twiddle_rsc_0_11_i_ARLEN <= twiddle_rsc_0_11_ARLEN;
  twiddle_rsc_0_11_i_ARSIZE <= twiddle_rsc_0_11_ARSIZE;
  twiddle_rsc_0_11_i_ARBURST <= twiddle_rsc_0_11_ARBURST;
  twiddle_rsc_0_11_i_ARCACHE <= twiddle_rsc_0_11_ARCACHE;
  twiddle_rsc_0_11_i_ARPROT <= twiddle_rsc_0_11_ARPROT;
  twiddle_rsc_0_11_i_ARQOS <= twiddle_rsc_0_11_ARQOS;
  twiddle_rsc_0_11_i_ARREGION <= twiddle_rsc_0_11_ARREGION;
  twiddle_rsc_0_11_i_ARUSER(0) <= twiddle_rsc_0_11_ARUSER;
  twiddle_rsc_0_11_RID <= twiddle_rsc_0_11_i_RID(0);
  twiddle_rsc_0_11_RDATA <= twiddle_rsc_0_11_i_RDATA;
  twiddle_rsc_0_11_RRESP <= twiddle_rsc_0_11_i_RRESP;
  twiddle_rsc_0_11_RUSER <= twiddle_rsc_0_11_i_RUSER(0);
  twiddle_rsc_0_11_i_s_raddr_1 <= twiddle_rsc_0_11_i_s_raddr;
  twiddle_rsc_0_11_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_11_i_s_din <= twiddle_rsc_0_11_i_s_din_1;
  twiddle_rsc_0_11_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_11_i_oswt => twiddle_rsc_0_11_i_oswt,
      twiddle_rsc_0_11_i_biwt => twiddle_rsc_0_11_i_biwt,
      twiddle_rsc_0_11_i_bdwt => twiddle_rsc_0_11_i_bdwt,
      twiddle_rsc_0_11_i_bcwt => twiddle_rsc_0_11_i_bcwt,
      twiddle_rsc_0_11_i_s_re_core_sct => twiddle_rsc_0_11_i_s_re_core_sct,
      twiddle_rsc_0_11_i_s_rrdy => twiddle_rsc_0_11_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_11_i_oswt => twiddle_rsc_0_11_i_oswt,
      twiddle_rsc_0_11_i_wen_comp => twiddle_rsc_0_11_i_wen_comp,
      twiddle_rsc_0_11_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp_inst_twiddle_rsc_0_11_i_s_raddr_core,
      twiddle_rsc_0_11_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp_inst_twiddle_rsc_0_11_i_s_din_mxwt,
      twiddle_rsc_0_11_i_biwt => twiddle_rsc_0_11_i_biwt,
      twiddle_rsc_0_11_i_bdwt => twiddle_rsc_0_11_i_bdwt,
      twiddle_rsc_0_11_i_bcwt => twiddle_rsc_0_11_i_bcwt,
      twiddle_rsc_0_11_i_s_raddr => peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp_inst_twiddle_rsc_0_11_i_s_raddr,
      twiddle_rsc_0_11_i_s_raddr_core_sct => twiddle_rsc_0_11_i_s_re_core_sct,
      twiddle_rsc_0_11_i_s_din => peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp_inst_twiddle_rsc_0_11_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp_inst_twiddle_rsc_0_11_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_11_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_11_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp_inst_twiddle_rsc_0_11_i_s_din_mxwt;
  twiddle_rsc_0_11_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp_inst_twiddle_rsc_0_11_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_11_i_twiddle_rsc_0_11_wait_dp_inst_twiddle_rsc_0_11_i_s_din
      <= twiddle_rsc_0_11_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_10_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_10_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_10_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_10_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_10_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_10_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_10_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_10_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_10_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_10_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_10_RID : OUT STD_LOGIC;
    twiddle_rsc_0_10_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_10_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_10_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_10_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_10_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_10_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_10_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_10_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_10_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_10_ARID : IN STD_LOGIC;
    twiddle_rsc_0_10_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_10_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_10_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_10_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_10_BID : OUT STD_LOGIC;
    twiddle_rsc_0_10_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_10_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_10_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_10_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_10_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_10_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_10_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_10_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_10_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_10_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_10_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_10_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_10_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_10_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_10_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_10_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_10_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_10_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_10_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_10_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_10_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_10_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_10_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_10_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_10_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_10_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_10_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_10_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_10_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_10_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_10_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_10_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_10_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_10_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_10_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_10_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_10_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_10_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_10_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_10_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_10_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_10_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_10_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_10_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_10_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp_inst_twiddle_rsc_0_10_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp_inst_twiddle_rsc_0_10_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp_inst_twiddle_rsc_0_10_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp_inst_twiddle_rsc_0_10_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_10_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_10_i_AWID,
      AWADDR => twiddle_rsc_0_10_i_AWADDR,
      AWLEN => twiddle_rsc_0_10_i_AWLEN,
      AWSIZE => twiddle_rsc_0_10_i_AWSIZE,
      AWBURST => twiddle_rsc_0_10_i_AWBURST,
      AWLOCK => twiddle_rsc_0_10_AWLOCK,
      AWCACHE => twiddle_rsc_0_10_i_AWCACHE,
      AWPROT => twiddle_rsc_0_10_i_AWPROT,
      AWQOS => twiddle_rsc_0_10_i_AWQOS,
      AWREGION => twiddle_rsc_0_10_i_AWREGION,
      AWUSER => twiddle_rsc_0_10_i_AWUSER,
      AWVALID => twiddle_rsc_0_10_AWVALID,
      AWREADY => twiddle_rsc_0_10_AWREADY,
      WDATA => twiddle_rsc_0_10_i_WDATA,
      WSTRB => twiddle_rsc_0_10_i_WSTRB,
      WLAST => twiddle_rsc_0_10_WLAST,
      WUSER => twiddle_rsc_0_10_i_WUSER,
      WVALID => twiddle_rsc_0_10_WVALID,
      WREADY => twiddle_rsc_0_10_WREADY,
      BID => twiddle_rsc_0_10_i_BID,
      BRESP => twiddle_rsc_0_10_i_BRESP,
      BUSER => twiddle_rsc_0_10_i_BUSER,
      BVALID => twiddle_rsc_0_10_BVALID,
      BREADY => twiddle_rsc_0_10_BREADY,
      ARID => twiddle_rsc_0_10_i_ARID,
      ARADDR => twiddle_rsc_0_10_i_ARADDR,
      ARLEN => twiddle_rsc_0_10_i_ARLEN,
      ARSIZE => twiddle_rsc_0_10_i_ARSIZE,
      ARBURST => twiddle_rsc_0_10_i_ARBURST,
      ARLOCK => twiddle_rsc_0_10_ARLOCK,
      ARCACHE => twiddle_rsc_0_10_i_ARCACHE,
      ARPROT => twiddle_rsc_0_10_i_ARPROT,
      ARQOS => twiddle_rsc_0_10_i_ARQOS,
      ARREGION => twiddle_rsc_0_10_i_ARREGION,
      ARUSER => twiddle_rsc_0_10_i_ARUSER,
      ARVALID => twiddle_rsc_0_10_ARVALID,
      ARREADY => twiddle_rsc_0_10_ARREADY,
      RID => twiddle_rsc_0_10_i_RID,
      RDATA => twiddle_rsc_0_10_i_RDATA,
      RRESP => twiddle_rsc_0_10_i_RRESP,
      RLAST => twiddle_rsc_0_10_RLAST,
      RUSER => twiddle_rsc_0_10_i_RUSER,
      RVALID => twiddle_rsc_0_10_RVALID,
      RREADY => twiddle_rsc_0_10_RREADY,
      s_re => twiddle_rsc_0_10_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_10_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_10_i_s_waddr,
      s_din => twiddle_rsc_0_10_i_s_din_1,
      s_dout => twiddle_rsc_0_10_i_s_dout,
      s_rrdy => twiddle_rsc_0_10_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_10_i_s_wrdy,
      is_idle => twiddle_rsc_0_10_is_idle,
      tr_write_done => twiddle_rsc_0_10_tr_write_done,
      s_tdone => twiddle_rsc_0_10_s_tdone
    );
  twiddle_rsc_0_10_i_AWID(0) <= twiddle_rsc_0_10_AWID;
  twiddle_rsc_0_10_i_AWADDR <= twiddle_rsc_0_10_AWADDR;
  twiddle_rsc_0_10_i_AWLEN <= twiddle_rsc_0_10_AWLEN;
  twiddle_rsc_0_10_i_AWSIZE <= twiddle_rsc_0_10_AWSIZE;
  twiddle_rsc_0_10_i_AWBURST <= twiddle_rsc_0_10_AWBURST;
  twiddle_rsc_0_10_i_AWCACHE <= twiddle_rsc_0_10_AWCACHE;
  twiddle_rsc_0_10_i_AWPROT <= twiddle_rsc_0_10_AWPROT;
  twiddle_rsc_0_10_i_AWQOS <= twiddle_rsc_0_10_AWQOS;
  twiddle_rsc_0_10_i_AWREGION <= twiddle_rsc_0_10_AWREGION;
  twiddle_rsc_0_10_i_AWUSER(0) <= twiddle_rsc_0_10_AWUSER;
  twiddle_rsc_0_10_i_WDATA <= twiddle_rsc_0_10_WDATA;
  twiddle_rsc_0_10_i_WSTRB <= twiddle_rsc_0_10_WSTRB;
  twiddle_rsc_0_10_i_WUSER(0) <= twiddle_rsc_0_10_WUSER;
  twiddle_rsc_0_10_BID <= twiddle_rsc_0_10_i_BID(0);
  twiddle_rsc_0_10_BRESP <= twiddle_rsc_0_10_i_BRESP;
  twiddle_rsc_0_10_BUSER <= twiddle_rsc_0_10_i_BUSER(0);
  twiddle_rsc_0_10_i_ARID(0) <= twiddle_rsc_0_10_ARID;
  twiddle_rsc_0_10_i_ARADDR <= twiddle_rsc_0_10_ARADDR;
  twiddle_rsc_0_10_i_ARLEN <= twiddle_rsc_0_10_ARLEN;
  twiddle_rsc_0_10_i_ARSIZE <= twiddle_rsc_0_10_ARSIZE;
  twiddle_rsc_0_10_i_ARBURST <= twiddle_rsc_0_10_ARBURST;
  twiddle_rsc_0_10_i_ARCACHE <= twiddle_rsc_0_10_ARCACHE;
  twiddle_rsc_0_10_i_ARPROT <= twiddle_rsc_0_10_ARPROT;
  twiddle_rsc_0_10_i_ARQOS <= twiddle_rsc_0_10_ARQOS;
  twiddle_rsc_0_10_i_ARREGION <= twiddle_rsc_0_10_ARREGION;
  twiddle_rsc_0_10_i_ARUSER(0) <= twiddle_rsc_0_10_ARUSER;
  twiddle_rsc_0_10_RID <= twiddle_rsc_0_10_i_RID(0);
  twiddle_rsc_0_10_RDATA <= twiddle_rsc_0_10_i_RDATA;
  twiddle_rsc_0_10_RRESP <= twiddle_rsc_0_10_i_RRESP;
  twiddle_rsc_0_10_RUSER <= twiddle_rsc_0_10_i_RUSER(0);
  twiddle_rsc_0_10_i_s_raddr_1 <= twiddle_rsc_0_10_i_s_raddr;
  twiddle_rsc_0_10_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_10_i_s_din <= twiddle_rsc_0_10_i_s_din_1;
  twiddle_rsc_0_10_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_10_i_oswt => twiddle_rsc_0_10_i_oswt,
      twiddle_rsc_0_10_i_biwt => twiddle_rsc_0_10_i_biwt,
      twiddle_rsc_0_10_i_bdwt => twiddle_rsc_0_10_i_bdwt,
      twiddle_rsc_0_10_i_bcwt => twiddle_rsc_0_10_i_bcwt,
      twiddle_rsc_0_10_i_s_re_core_sct => twiddle_rsc_0_10_i_s_re_core_sct,
      twiddle_rsc_0_10_i_s_rrdy => twiddle_rsc_0_10_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_10_i_oswt => twiddle_rsc_0_10_i_oswt,
      twiddle_rsc_0_10_i_wen_comp => twiddle_rsc_0_10_i_wen_comp,
      twiddle_rsc_0_10_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp_inst_twiddle_rsc_0_10_i_s_raddr_core,
      twiddle_rsc_0_10_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp_inst_twiddle_rsc_0_10_i_s_din_mxwt,
      twiddle_rsc_0_10_i_biwt => twiddle_rsc_0_10_i_biwt,
      twiddle_rsc_0_10_i_bdwt => twiddle_rsc_0_10_i_bdwt,
      twiddle_rsc_0_10_i_bcwt => twiddle_rsc_0_10_i_bcwt,
      twiddle_rsc_0_10_i_s_raddr => peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp_inst_twiddle_rsc_0_10_i_s_raddr,
      twiddle_rsc_0_10_i_s_raddr_core_sct => twiddle_rsc_0_10_i_s_re_core_sct,
      twiddle_rsc_0_10_i_s_din => peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp_inst_twiddle_rsc_0_10_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp_inst_twiddle_rsc_0_10_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_10_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_10_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp_inst_twiddle_rsc_0_10_i_s_din_mxwt;
  twiddle_rsc_0_10_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp_inst_twiddle_rsc_0_10_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_10_i_twiddle_rsc_0_10_wait_dp_inst_twiddle_rsc_0_10_i_s_din
      <= twiddle_rsc_0_10_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_9_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_9_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_9_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_9_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_9_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_9_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_9_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_9_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_9_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_9_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_9_RID : OUT STD_LOGIC;
    twiddle_rsc_0_9_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_9_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_9_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_9_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_9_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_9_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_9_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_9_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_9_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_9_ARID : IN STD_LOGIC;
    twiddle_rsc_0_9_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_9_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_9_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_9_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_9_BID : OUT STD_LOGIC;
    twiddle_rsc_0_9_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_9_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_9_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_9_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_9_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_9_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_9_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_9_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_9_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_9_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_9_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_9_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_9_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_9_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_9_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_9_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_9_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_9_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_9_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_9_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_9_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_9_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_9_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_9_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_9_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_9_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_9_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_9_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_9_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_9_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_9_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_9_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_9_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_9_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_9_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_9_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_9_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_9_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_9_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_9_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_9_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_9_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_9_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_9_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_9_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp_inst_twiddle_rsc_0_9_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp_inst_twiddle_rsc_0_9_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp_inst_twiddle_rsc_0_9_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp_inst_twiddle_rsc_0_9_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_9_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_9_i_AWID,
      AWADDR => twiddle_rsc_0_9_i_AWADDR,
      AWLEN => twiddle_rsc_0_9_i_AWLEN,
      AWSIZE => twiddle_rsc_0_9_i_AWSIZE,
      AWBURST => twiddle_rsc_0_9_i_AWBURST,
      AWLOCK => twiddle_rsc_0_9_AWLOCK,
      AWCACHE => twiddle_rsc_0_9_i_AWCACHE,
      AWPROT => twiddle_rsc_0_9_i_AWPROT,
      AWQOS => twiddle_rsc_0_9_i_AWQOS,
      AWREGION => twiddle_rsc_0_9_i_AWREGION,
      AWUSER => twiddle_rsc_0_9_i_AWUSER,
      AWVALID => twiddle_rsc_0_9_AWVALID,
      AWREADY => twiddle_rsc_0_9_AWREADY,
      WDATA => twiddle_rsc_0_9_i_WDATA,
      WSTRB => twiddle_rsc_0_9_i_WSTRB,
      WLAST => twiddle_rsc_0_9_WLAST,
      WUSER => twiddle_rsc_0_9_i_WUSER,
      WVALID => twiddle_rsc_0_9_WVALID,
      WREADY => twiddle_rsc_0_9_WREADY,
      BID => twiddle_rsc_0_9_i_BID,
      BRESP => twiddle_rsc_0_9_i_BRESP,
      BUSER => twiddle_rsc_0_9_i_BUSER,
      BVALID => twiddle_rsc_0_9_BVALID,
      BREADY => twiddle_rsc_0_9_BREADY,
      ARID => twiddle_rsc_0_9_i_ARID,
      ARADDR => twiddle_rsc_0_9_i_ARADDR,
      ARLEN => twiddle_rsc_0_9_i_ARLEN,
      ARSIZE => twiddle_rsc_0_9_i_ARSIZE,
      ARBURST => twiddle_rsc_0_9_i_ARBURST,
      ARLOCK => twiddle_rsc_0_9_ARLOCK,
      ARCACHE => twiddle_rsc_0_9_i_ARCACHE,
      ARPROT => twiddle_rsc_0_9_i_ARPROT,
      ARQOS => twiddle_rsc_0_9_i_ARQOS,
      ARREGION => twiddle_rsc_0_9_i_ARREGION,
      ARUSER => twiddle_rsc_0_9_i_ARUSER,
      ARVALID => twiddle_rsc_0_9_ARVALID,
      ARREADY => twiddle_rsc_0_9_ARREADY,
      RID => twiddle_rsc_0_9_i_RID,
      RDATA => twiddle_rsc_0_9_i_RDATA,
      RRESP => twiddle_rsc_0_9_i_RRESP,
      RLAST => twiddle_rsc_0_9_RLAST,
      RUSER => twiddle_rsc_0_9_i_RUSER,
      RVALID => twiddle_rsc_0_9_RVALID,
      RREADY => twiddle_rsc_0_9_RREADY,
      s_re => twiddle_rsc_0_9_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_9_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_9_i_s_waddr,
      s_din => twiddle_rsc_0_9_i_s_din_1,
      s_dout => twiddle_rsc_0_9_i_s_dout,
      s_rrdy => twiddle_rsc_0_9_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_9_i_s_wrdy,
      is_idle => twiddle_rsc_0_9_is_idle,
      tr_write_done => twiddle_rsc_0_9_tr_write_done,
      s_tdone => twiddle_rsc_0_9_s_tdone
    );
  twiddle_rsc_0_9_i_AWID(0) <= twiddle_rsc_0_9_AWID;
  twiddle_rsc_0_9_i_AWADDR <= twiddle_rsc_0_9_AWADDR;
  twiddle_rsc_0_9_i_AWLEN <= twiddle_rsc_0_9_AWLEN;
  twiddle_rsc_0_9_i_AWSIZE <= twiddle_rsc_0_9_AWSIZE;
  twiddle_rsc_0_9_i_AWBURST <= twiddle_rsc_0_9_AWBURST;
  twiddle_rsc_0_9_i_AWCACHE <= twiddle_rsc_0_9_AWCACHE;
  twiddle_rsc_0_9_i_AWPROT <= twiddle_rsc_0_9_AWPROT;
  twiddle_rsc_0_9_i_AWQOS <= twiddle_rsc_0_9_AWQOS;
  twiddle_rsc_0_9_i_AWREGION <= twiddle_rsc_0_9_AWREGION;
  twiddle_rsc_0_9_i_AWUSER(0) <= twiddle_rsc_0_9_AWUSER;
  twiddle_rsc_0_9_i_WDATA <= twiddle_rsc_0_9_WDATA;
  twiddle_rsc_0_9_i_WSTRB <= twiddle_rsc_0_9_WSTRB;
  twiddle_rsc_0_9_i_WUSER(0) <= twiddle_rsc_0_9_WUSER;
  twiddle_rsc_0_9_BID <= twiddle_rsc_0_9_i_BID(0);
  twiddle_rsc_0_9_BRESP <= twiddle_rsc_0_9_i_BRESP;
  twiddle_rsc_0_9_BUSER <= twiddle_rsc_0_9_i_BUSER(0);
  twiddle_rsc_0_9_i_ARID(0) <= twiddle_rsc_0_9_ARID;
  twiddle_rsc_0_9_i_ARADDR <= twiddle_rsc_0_9_ARADDR;
  twiddle_rsc_0_9_i_ARLEN <= twiddle_rsc_0_9_ARLEN;
  twiddle_rsc_0_9_i_ARSIZE <= twiddle_rsc_0_9_ARSIZE;
  twiddle_rsc_0_9_i_ARBURST <= twiddle_rsc_0_9_ARBURST;
  twiddle_rsc_0_9_i_ARCACHE <= twiddle_rsc_0_9_ARCACHE;
  twiddle_rsc_0_9_i_ARPROT <= twiddle_rsc_0_9_ARPROT;
  twiddle_rsc_0_9_i_ARQOS <= twiddle_rsc_0_9_ARQOS;
  twiddle_rsc_0_9_i_ARREGION <= twiddle_rsc_0_9_ARREGION;
  twiddle_rsc_0_9_i_ARUSER(0) <= twiddle_rsc_0_9_ARUSER;
  twiddle_rsc_0_9_RID <= twiddle_rsc_0_9_i_RID(0);
  twiddle_rsc_0_9_RDATA <= twiddle_rsc_0_9_i_RDATA;
  twiddle_rsc_0_9_RRESP <= twiddle_rsc_0_9_i_RRESP;
  twiddle_rsc_0_9_RUSER <= twiddle_rsc_0_9_i_RUSER(0);
  twiddle_rsc_0_9_i_s_raddr_1 <= twiddle_rsc_0_9_i_s_raddr;
  twiddle_rsc_0_9_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_9_i_s_din <= twiddle_rsc_0_9_i_s_din_1;
  twiddle_rsc_0_9_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_9_i_oswt => twiddle_rsc_0_9_i_oswt,
      twiddle_rsc_0_9_i_biwt => twiddle_rsc_0_9_i_biwt,
      twiddle_rsc_0_9_i_bdwt => twiddle_rsc_0_9_i_bdwt,
      twiddle_rsc_0_9_i_bcwt => twiddle_rsc_0_9_i_bcwt,
      twiddle_rsc_0_9_i_s_re_core_sct => twiddle_rsc_0_9_i_s_re_core_sct,
      twiddle_rsc_0_9_i_s_rrdy => twiddle_rsc_0_9_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_9_i_oswt => twiddle_rsc_0_9_i_oswt,
      twiddle_rsc_0_9_i_wen_comp => twiddle_rsc_0_9_i_wen_comp,
      twiddle_rsc_0_9_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp_inst_twiddle_rsc_0_9_i_s_raddr_core,
      twiddle_rsc_0_9_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp_inst_twiddle_rsc_0_9_i_s_din_mxwt,
      twiddle_rsc_0_9_i_biwt => twiddle_rsc_0_9_i_biwt,
      twiddle_rsc_0_9_i_bdwt => twiddle_rsc_0_9_i_bdwt,
      twiddle_rsc_0_9_i_bcwt => twiddle_rsc_0_9_i_bcwt,
      twiddle_rsc_0_9_i_s_raddr => peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp_inst_twiddle_rsc_0_9_i_s_raddr,
      twiddle_rsc_0_9_i_s_raddr_core_sct => twiddle_rsc_0_9_i_s_re_core_sct,
      twiddle_rsc_0_9_i_s_din => peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp_inst_twiddle_rsc_0_9_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp_inst_twiddle_rsc_0_9_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_9_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_9_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp_inst_twiddle_rsc_0_9_i_s_din_mxwt;
  twiddle_rsc_0_9_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp_inst_twiddle_rsc_0_9_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_9_i_twiddle_rsc_0_9_wait_dp_inst_twiddle_rsc_0_9_i_s_din
      <= twiddle_rsc_0_9_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_8_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_8_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_8_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_8_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_8_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_8_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_8_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_8_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_8_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_8_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_8_RID : OUT STD_LOGIC;
    twiddle_rsc_0_8_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_8_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_8_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_8_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_8_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_8_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_8_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_8_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_8_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_8_ARID : IN STD_LOGIC;
    twiddle_rsc_0_8_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_8_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_8_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_8_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_8_BID : OUT STD_LOGIC;
    twiddle_rsc_0_8_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_8_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_8_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_8_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_8_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_8_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_8_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_8_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_8_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_8_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_8_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_8_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_8_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_8_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_8_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_8_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_8_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_8_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_8_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_8_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_8_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_8_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_8_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_8_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_8_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_8_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_8_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_8_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_8_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_8_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_8_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_8_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_8_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_8_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_8_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_8_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_8_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_8_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_8_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_8_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_8_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_8_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_8_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_8_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_8_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp_inst_twiddle_rsc_0_8_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp_inst_twiddle_rsc_0_8_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp_inst_twiddle_rsc_0_8_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp_inst_twiddle_rsc_0_8_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_8_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_8_i_AWID,
      AWADDR => twiddle_rsc_0_8_i_AWADDR,
      AWLEN => twiddle_rsc_0_8_i_AWLEN,
      AWSIZE => twiddle_rsc_0_8_i_AWSIZE,
      AWBURST => twiddle_rsc_0_8_i_AWBURST,
      AWLOCK => twiddle_rsc_0_8_AWLOCK,
      AWCACHE => twiddle_rsc_0_8_i_AWCACHE,
      AWPROT => twiddle_rsc_0_8_i_AWPROT,
      AWQOS => twiddle_rsc_0_8_i_AWQOS,
      AWREGION => twiddle_rsc_0_8_i_AWREGION,
      AWUSER => twiddle_rsc_0_8_i_AWUSER,
      AWVALID => twiddle_rsc_0_8_AWVALID,
      AWREADY => twiddle_rsc_0_8_AWREADY,
      WDATA => twiddle_rsc_0_8_i_WDATA,
      WSTRB => twiddle_rsc_0_8_i_WSTRB,
      WLAST => twiddle_rsc_0_8_WLAST,
      WUSER => twiddle_rsc_0_8_i_WUSER,
      WVALID => twiddle_rsc_0_8_WVALID,
      WREADY => twiddle_rsc_0_8_WREADY,
      BID => twiddle_rsc_0_8_i_BID,
      BRESP => twiddle_rsc_0_8_i_BRESP,
      BUSER => twiddle_rsc_0_8_i_BUSER,
      BVALID => twiddle_rsc_0_8_BVALID,
      BREADY => twiddle_rsc_0_8_BREADY,
      ARID => twiddle_rsc_0_8_i_ARID,
      ARADDR => twiddle_rsc_0_8_i_ARADDR,
      ARLEN => twiddle_rsc_0_8_i_ARLEN,
      ARSIZE => twiddle_rsc_0_8_i_ARSIZE,
      ARBURST => twiddle_rsc_0_8_i_ARBURST,
      ARLOCK => twiddle_rsc_0_8_ARLOCK,
      ARCACHE => twiddle_rsc_0_8_i_ARCACHE,
      ARPROT => twiddle_rsc_0_8_i_ARPROT,
      ARQOS => twiddle_rsc_0_8_i_ARQOS,
      ARREGION => twiddle_rsc_0_8_i_ARREGION,
      ARUSER => twiddle_rsc_0_8_i_ARUSER,
      ARVALID => twiddle_rsc_0_8_ARVALID,
      ARREADY => twiddle_rsc_0_8_ARREADY,
      RID => twiddle_rsc_0_8_i_RID,
      RDATA => twiddle_rsc_0_8_i_RDATA,
      RRESP => twiddle_rsc_0_8_i_RRESP,
      RLAST => twiddle_rsc_0_8_RLAST,
      RUSER => twiddle_rsc_0_8_i_RUSER,
      RVALID => twiddle_rsc_0_8_RVALID,
      RREADY => twiddle_rsc_0_8_RREADY,
      s_re => twiddle_rsc_0_8_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_8_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_8_i_s_waddr,
      s_din => twiddle_rsc_0_8_i_s_din_1,
      s_dout => twiddle_rsc_0_8_i_s_dout,
      s_rrdy => twiddle_rsc_0_8_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_8_i_s_wrdy,
      is_idle => twiddle_rsc_0_8_is_idle,
      tr_write_done => twiddle_rsc_0_8_tr_write_done,
      s_tdone => twiddle_rsc_0_8_s_tdone
    );
  twiddle_rsc_0_8_i_AWID(0) <= twiddle_rsc_0_8_AWID;
  twiddle_rsc_0_8_i_AWADDR <= twiddle_rsc_0_8_AWADDR;
  twiddle_rsc_0_8_i_AWLEN <= twiddle_rsc_0_8_AWLEN;
  twiddle_rsc_0_8_i_AWSIZE <= twiddle_rsc_0_8_AWSIZE;
  twiddle_rsc_0_8_i_AWBURST <= twiddle_rsc_0_8_AWBURST;
  twiddle_rsc_0_8_i_AWCACHE <= twiddle_rsc_0_8_AWCACHE;
  twiddle_rsc_0_8_i_AWPROT <= twiddle_rsc_0_8_AWPROT;
  twiddle_rsc_0_8_i_AWQOS <= twiddle_rsc_0_8_AWQOS;
  twiddle_rsc_0_8_i_AWREGION <= twiddle_rsc_0_8_AWREGION;
  twiddle_rsc_0_8_i_AWUSER(0) <= twiddle_rsc_0_8_AWUSER;
  twiddle_rsc_0_8_i_WDATA <= twiddle_rsc_0_8_WDATA;
  twiddle_rsc_0_8_i_WSTRB <= twiddle_rsc_0_8_WSTRB;
  twiddle_rsc_0_8_i_WUSER(0) <= twiddle_rsc_0_8_WUSER;
  twiddle_rsc_0_8_BID <= twiddle_rsc_0_8_i_BID(0);
  twiddle_rsc_0_8_BRESP <= twiddle_rsc_0_8_i_BRESP;
  twiddle_rsc_0_8_BUSER <= twiddle_rsc_0_8_i_BUSER(0);
  twiddle_rsc_0_8_i_ARID(0) <= twiddle_rsc_0_8_ARID;
  twiddle_rsc_0_8_i_ARADDR <= twiddle_rsc_0_8_ARADDR;
  twiddle_rsc_0_8_i_ARLEN <= twiddle_rsc_0_8_ARLEN;
  twiddle_rsc_0_8_i_ARSIZE <= twiddle_rsc_0_8_ARSIZE;
  twiddle_rsc_0_8_i_ARBURST <= twiddle_rsc_0_8_ARBURST;
  twiddle_rsc_0_8_i_ARCACHE <= twiddle_rsc_0_8_ARCACHE;
  twiddle_rsc_0_8_i_ARPROT <= twiddle_rsc_0_8_ARPROT;
  twiddle_rsc_0_8_i_ARQOS <= twiddle_rsc_0_8_ARQOS;
  twiddle_rsc_0_8_i_ARREGION <= twiddle_rsc_0_8_ARREGION;
  twiddle_rsc_0_8_i_ARUSER(0) <= twiddle_rsc_0_8_ARUSER;
  twiddle_rsc_0_8_RID <= twiddle_rsc_0_8_i_RID(0);
  twiddle_rsc_0_8_RDATA <= twiddle_rsc_0_8_i_RDATA;
  twiddle_rsc_0_8_RRESP <= twiddle_rsc_0_8_i_RRESP;
  twiddle_rsc_0_8_RUSER <= twiddle_rsc_0_8_i_RUSER(0);
  twiddle_rsc_0_8_i_s_raddr_1 <= twiddle_rsc_0_8_i_s_raddr;
  twiddle_rsc_0_8_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_8_i_s_din <= twiddle_rsc_0_8_i_s_din_1;
  twiddle_rsc_0_8_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_8_i_oswt => twiddle_rsc_0_8_i_oswt,
      twiddle_rsc_0_8_i_biwt => twiddle_rsc_0_8_i_biwt,
      twiddle_rsc_0_8_i_bdwt => twiddle_rsc_0_8_i_bdwt,
      twiddle_rsc_0_8_i_bcwt => twiddle_rsc_0_8_i_bcwt,
      twiddle_rsc_0_8_i_s_re_core_sct => twiddle_rsc_0_8_i_s_re_core_sct,
      twiddle_rsc_0_8_i_s_rrdy => twiddle_rsc_0_8_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_8_i_oswt => twiddle_rsc_0_8_i_oswt,
      twiddle_rsc_0_8_i_wen_comp => twiddle_rsc_0_8_i_wen_comp,
      twiddle_rsc_0_8_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp_inst_twiddle_rsc_0_8_i_s_raddr_core,
      twiddle_rsc_0_8_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp_inst_twiddle_rsc_0_8_i_s_din_mxwt,
      twiddle_rsc_0_8_i_biwt => twiddle_rsc_0_8_i_biwt,
      twiddle_rsc_0_8_i_bdwt => twiddle_rsc_0_8_i_bdwt,
      twiddle_rsc_0_8_i_bcwt => twiddle_rsc_0_8_i_bcwt,
      twiddle_rsc_0_8_i_s_raddr => peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp_inst_twiddle_rsc_0_8_i_s_raddr,
      twiddle_rsc_0_8_i_s_raddr_core_sct => twiddle_rsc_0_8_i_s_re_core_sct,
      twiddle_rsc_0_8_i_s_din => peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp_inst_twiddle_rsc_0_8_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp_inst_twiddle_rsc_0_8_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_8_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_8_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp_inst_twiddle_rsc_0_8_i_s_din_mxwt;
  twiddle_rsc_0_8_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp_inst_twiddle_rsc_0_8_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_8_i_twiddle_rsc_0_8_wait_dp_inst_twiddle_rsc_0_8_i_s_din
      <= twiddle_rsc_0_8_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_7_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_7_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_7_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_7_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_7_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_7_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_7_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_7_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_7_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_7_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_RID : OUT STD_LOGIC;
    twiddle_rsc_0_7_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_7_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_7_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_7_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_7_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_7_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_7_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_7_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_7_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_7_ARID : IN STD_LOGIC;
    twiddle_rsc_0_7_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_7_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_7_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_7_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_7_BID : OUT STD_LOGIC;
    twiddle_rsc_0_7_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_7_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_7_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_7_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_7_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_7_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_7_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_7_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_7_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_7_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_7_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_7_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_7_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_7_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_7_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_7_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_7_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_7_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_7_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_7_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_7_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_7_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_7_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_7_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_7_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_7_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_7_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_7_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_7_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_7_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_7_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_7_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_7_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_7_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_7_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_7_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_7_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_7_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_7_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_7_i_AWID,
      AWADDR => twiddle_rsc_0_7_i_AWADDR,
      AWLEN => twiddle_rsc_0_7_i_AWLEN,
      AWSIZE => twiddle_rsc_0_7_i_AWSIZE,
      AWBURST => twiddle_rsc_0_7_i_AWBURST,
      AWLOCK => twiddle_rsc_0_7_AWLOCK,
      AWCACHE => twiddle_rsc_0_7_i_AWCACHE,
      AWPROT => twiddle_rsc_0_7_i_AWPROT,
      AWQOS => twiddle_rsc_0_7_i_AWQOS,
      AWREGION => twiddle_rsc_0_7_i_AWREGION,
      AWUSER => twiddle_rsc_0_7_i_AWUSER,
      AWVALID => twiddle_rsc_0_7_AWVALID,
      AWREADY => twiddle_rsc_0_7_AWREADY,
      WDATA => twiddle_rsc_0_7_i_WDATA,
      WSTRB => twiddle_rsc_0_7_i_WSTRB,
      WLAST => twiddle_rsc_0_7_WLAST,
      WUSER => twiddle_rsc_0_7_i_WUSER,
      WVALID => twiddle_rsc_0_7_WVALID,
      WREADY => twiddle_rsc_0_7_WREADY,
      BID => twiddle_rsc_0_7_i_BID,
      BRESP => twiddle_rsc_0_7_i_BRESP,
      BUSER => twiddle_rsc_0_7_i_BUSER,
      BVALID => twiddle_rsc_0_7_BVALID,
      BREADY => twiddle_rsc_0_7_BREADY,
      ARID => twiddle_rsc_0_7_i_ARID,
      ARADDR => twiddle_rsc_0_7_i_ARADDR,
      ARLEN => twiddle_rsc_0_7_i_ARLEN,
      ARSIZE => twiddle_rsc_0_7_i_ARSIZE,
      ARBURST => twiddle_rsc_0_7_i_ARBURST,
      ARLOCK => twiddle_rsc_0_7_ARLOCK,
      ARCACHE => twiddle_rsc_0_7_i_ARCACHE,
      ARPROT => twiddle_rsc_0_7_i_ARPROT,
      ARQOS => twiddle_rsc_0_7_i_ARQOS,
      ARREGION => twiddle_rsc_0_7_i_ARREGION,
      ARUSER => twiddle_rsc_0_7_i_ARUSER,
      ARVALID => twiddle_rsc_0_7_ARVALID,
      ARREADY => twiddle_rsc_0_7_ARREADY,
      RID => twiddle_rsc_0_7_i_RID,
      RDATA => twiddle_rsc_0_7_i_RDATA,
      RRESP => twiddle_rsc_0_7_i_RRESP,
      RLAST => twiddle_rsc_0_7_RLAST,
      RUSER => twiddle_rsc_0_7_i_RUSER,
      RVALID => twiddle_rsc_0_7_RVALID,
      RREADY => twiddle_rsc_0_7_RREADY,
      s_re => twiddle_rsc_0_7_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_7_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_7_i_s_waddr,
      s_din => twiddle_rsc_0_7_i_s_din_1,
      s_dout => twiddle_rsc_0_7_i_s_dout,
      s_rrdy => twiddle_rsc_0_7_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_7_i_s_wrdy,
      is_idle => twiddle_rsc_0_7_is_idle,
      tr_write_done => twiddle_rsc_0_7_tr_write_done,
      s_tdone => twiddle_rsc_0_7_s_tdone
    );
  twiddle_rsc_0_7_i_AWID(0) <= twiddle_rsc_0_7_AWID;
  twiddle_rsc_0_7_i_AWADDR <= twiddle_rsc_0_7_AWADDR;
  twiddle_rsc_0_7_i_AWLEN <= twiddle_rsc_0_7_AWLEN;
  twiddle_rsc_0_7_i_AWSIZE <= twiddle_rsc_0_7_AWSIZE;
  twiddle_rsc_0_7_i_AWBURST <= twiddle_rsc_0_7_AWBURST;
  twiddle_rsc_0_7_i_AWCACHE <= twiddle_rsc_0_7_AWCACHE;
  twiddle_rsc_0_7_i_AWPROT <= twiddle_rsc_0_7_AWPROT;
  twiddle_rsc_0_7_i_AWQOS <= twiddle_rsc_0_7_AWQOS;
  twiddle_rsc_0_7_i_AWREGION <= twiddle_rsc_0_7_AWREGION;
  twiddle_rsc_0_7_i_AWUSER(0) <= twiddle_rsc_0_7_AWUSER;
  twiddle_rsc_0_7_i_WDATA <= twiddle_rsc_0_7_WDATA;
  twiddle_rsc_0_7_i_WSTRB <= twiddle_rsc_0_7_WSTRB;
  twiddle_rsc_0_7_i_WUSER(0) <= twiddle_rsc_0_7_WUSER;
  twiddle_rsc_0_7_BID <= twiddle_rsc_0_7_i_BID(0);
  twiddle_rsc_0_7_BRESP <= twiddle_rsc_0_7_i_BRESP;
  twiddle_rsc_0_7_BUSER <= twiddle_rsc_0_7_i_BUSER(0);
  twiddle_rsc_0_7_i_ARID(0) <= twiddle_rsc_0_7_ARID;
  twiddle_rsc_0_7_i_ARADDR <= twiddle_rsc_0_7_ARADDR;
  twiddle_rsc_0_7_i_ARLEN <= twiddle_rsc_0_7_ARLEN;
  twiddle_rsc_0_7_i_ARSIZE <= twiddle_rsc_0_7_ARSIZE;
  twiddle_rsc_0_7_i_ARBURST <= twiddle_rsc_0_7_ARBURST;
  twiddle_rsc_0_7_i_ARCACHE <= twiddle_rsc_0_7_ARCACHE;
  twiddle_rsc_0_7_i_ARPROT <= twiddle_rsc_0_7_ARPROT;
  twiddle_rsc_0_7_i_ARQOS <= twiddle_rsc_0_7_ARQOS;
  twiddle_rsc_0_7_i_ARREGION <= twiddle_rsc_0_7_ARREGION;
  twiddle_rsc_0_7_i_ARUSER(0) <= twiddle_rsc_0_7_ARUSER;
  twiddle_rsc_0_7_RID <= twiddle_rsc_0_7_i_RID(0);
  twiddle_rsc_0_7_RDATA <= twiddle_rsc_0_7_i_RDATA;
  twiddle_rsc_0_7_RRESP <= twiddle_rsc_0_7_i_RRESP;
  twiddle_rsc_0_7_RUSER <= twiddle_rsc_0_7_i_RUSER(0);
  twiddle_rsc_0_7_i_s_raddr_1 <= twiddle_rsc_0_7_i_s_raddr;
  twiddle_rsc_0_7_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_7_i_s_din <= twiddle_rsc_0_7_i_s_din_1;
  twiddle_rsc_0_7_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_7_i_oswt => twiddle_rsc_0_7_i_oswt,
      twiddle_rsc_0_7_i_biwt => twiddle_rsc_0_7_i_biwt,
      twiddle_rsc_0_7_i_bdwt => twiddle_rsc_0_7_i_bdwt,
      twiddle_rsc_0_7_i_bcwt => twiddle_rsc_0_7_i_bcwt,
      twiddle_rsc_0_7_i_s_re_core_sct => twiddle_rsc_0_7_i_s_re_core_sct,
      twiddle_rsc_0_7_i_s_rrdy => twiddle_rsc_0_7_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_7_i_oswt => twiddle_rsc_0_7_i_oswt,
      twiddle_rsc_0_7_i_wen_comp => twiddle_rsc_0_7_i_wen_comp,
      twiddle_rsc_0_7_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_s_raddr_core,
      twiddle_rsc_0_7_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_s_din_mxwt,
      twiddle_rsc_0_7_i_biwt => twiddle_rsc_0_7_i_biwt,
      twiddle_rsc_0_7_i_bdwt => twiddle_rsc_0_7_i_bdwt,
      twiddle_rsc_0_7_i_bcwt => twiddle_rsc_0_7_i_bcwt,
      twiddle_rsc_0_7_i_s_raddr => peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_s_raddr,
      twiddle_rsc_0_7_i_s_raddr_core_sct => twiddle_rsc_0_7_i_s_re_core_sct,
      twiddle_rsc_0_7_i_s_din => peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_7_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_7_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_s_din_mxwt;
  twiddle_rsc_0_7_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_7_i_twiddle_rsc_0_7_wait_dp_inst_twiddle_rsc_0_7_i_s_din
      <= twiddle_rsc_0_7_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_6_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_6_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_6_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_6_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_6_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_6_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_6_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_6_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_6_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_6_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_RID : OUT STD_LOGIC;
    twiddle_rsc_0_6_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_6_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_6_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_6_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_6_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_6_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_6_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_6_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_6_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_6_ARID : IN STD_LOGIC;
    twiddle_rsc_0_6_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_6_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_6_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_6_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_6_BID : OUT STD_LOGIC;
    twiddle_rsc_0_6_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_6_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_6_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_6_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_6_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_6_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_6_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_6_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_6_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_6_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_6_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_6_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_6_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_6_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_6_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_6_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_6_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_6_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_6_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_6_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_6_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_6_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_6_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_6_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_6_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_6_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_6_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_6_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_6_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_6_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_6_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_6_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_6_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_6_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_6_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_6_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_6_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_6_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_6_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_6_i_AWID,
      AWADDR => twiddle_rsc_0_6_i_AWADDR,
      AWLEN => twiddle_rsc_0_6_i_AWLEN,
      AWSIZE => twiddle_rsc_0_6_i_AWSIZE,
      AWBURST => twiddle_rsc_0_6_i_AWBURST,
      AWLOCK => twiddle_rsc_0_6_AWLOCK,
      AWCACHE => twiddle_rsc_0_6_i_AWCACHE,
      AWPROT => twiddle_rsc_0_6_i_AWPROT,
      AWQOS => twiddle_rsc_0_6_i_AWQOS,
      AWREGION => twiddle_rsc_0_6_i_AWREGION,
      AWUSER => twiddle_rsc_0_6_i_AWUSER,
      AWVALID => twiddle_rsc_0_6_AWVALID,
      AWREADY => twiddle_rsc_0_6_AWREADY,
      WDATA => twiddle_rsc_0_6_i_WDATA,
      WSTRB => twiddle_rsc_0_6_i_WSTRB,
      WLAST => twiddle_rsc_0_6_WLAST,
      WUSER => twiddle_rsc_0_6_i_WUSER,
      WVALID => twiddle_rsc_0_6_WVALID,
      WREADY => twiddle_rsc_0_6_WREADY,
      BID => twiddle_rsc_0_6_i_BID,
      BRESP => twiddle_rsc_0_6_i_BRESP,
      BUSER => twiddle_rsc_0_6_i_BUSER,
      BVALID => twiddle_rsc_0_6_BVALID,
      BREADY => twiddle_rsc_0_6_BREADY,
      ARID => twiddle_rsc_0_6_i_ARID,
      ARADDR => twiddle_rsc_0_6_i_ARADDR,
      ARLEN => twiddle_rsc_0_6_i_ARLEN,
      ARSIZE => twiddle_rsc_0_6_i_ARSIZE,
      ARBURST => twiddle_rsc_0_6_i_ARBURST,
      ARLOCK => twiddle_rsc_0_6_ARLOCK,
      ARCACHE => twiddle_rsc_0_6_i_ARCACHE,
      ARPROT => twiddle_rsc_0_6_i_ARPROT,
      ARQOS => twiddle_rsc_0_6_i_ARQOS,
      ARREGION => twiddle_rsc_0_6_i_ARREGION,
      ARUSER => twiddle_rsc_0_6_i_ARUSER,
      ARVALID => twiddle_rsc_0_6_ARVALID,
      ARREADY => twiddle_rsc_0_6_ARREADY,
      RID => twiddle_rsc_0_6_i_RID,
      RDATA => twiddle_rsc_0_6_i_RDATA,
      RRESP => twiddle_rsc_0_6_i_RRESP,
      RLAST => twiddle_rsc_0_6_RLAST,
      RUSER => twiddle_rsc_0_6_i_RUSER,
      RVALID => twiddle_rsc_0_6_RVALID,
      RREADY => twiddle_rsc_0_6_RREADY,
      s_re => twiddle_rsc_0_6_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_6_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_6_i_s_waddr,
      s_din => twiddle_rsc_0_6_i_s_din_1,
      s_dout => twiddle_rsc_0_6_i_s_dout,
      s_rrdy => twiddle_rsc_0_6_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_6_i_s_wrdy,
      is_idle => twiddle_rsc_0_6_is_idle,
      tr_write_done => twiddle_rsc_0_6_tr_write_done,
      s_tdone => twiddle_rsc_0_6_s_tdone
    );
  twiddle_rsc_0_6_i_AWID(0) <= twiddle_rsc_0_6_AWID;
  twiddle_rsc_0_6_i_AWADDR <= twiddle_rsc_0_6_AWADDR;
  twiddle_rsc_0_6_i_AWLEN <= twiddle_rsc_0_6_AWLEN;
  twiddle_rsc_0_6_i_AWSIZE <= twiddle_rsc_0_6_AWSIZE;
  twiddle_rsc_0_6_i_AWBURST <= twiddle_rsc_0_6_AWBURST;
  twiddle_rsc_0_6_i_AWCACHE <= twiddle_rsc_0_6_AWCACHE;
  twiddle_rsc_0_6_i_AWPROT <= twiddle_rsc_0_6_AWPROT;
  twiddle_rsc_0_6_i_AWQOS <= twiddle_rsc_0_6_AWQOS;
  twiddle_rsc_0_6_i_AWREGION <= twiddle_rsc_0_6_AWREGION;
  twiddle_rsc_0_6_i_AWUSER(0) <= twiddle_rsc_0_6_AWUSER;
  twiddle_rsc_0_6_i_WDATA <= twiddle_rsc_0_6_WDATA;
  twiddle_rsc_0_6_i_WSTRB <= twiddle_rsc_0_6_WSTRB;
  twiddle_rsc_0_6_i_WUSER(0) <= twiddle_rsc_0_6_WUSER;
  twiddle_rsc_0_6_BID <= twiddle_rsc_0_6_i_BID(0);
  twiddle_rsc_0_6_BRESP <= twiddle_rsc_0_6_i_BRESP;
  twiddle_rsc_0_6_BUSER <= twiddle_rsc_0_6_i_BUSER(0);
  twiddle_rsc_0_6_i_ARID(0) <= twiddle_rsc_0_6_ARID;
  twiddle_rsc_0_6_i_ARADDR <= twiddle_rsc_0_6_ARADDR;
  twiddle_rsc_0_6_i_ARLEN <= twiddle_rsc_0_6_ARLEN;
  twiddle_rsc_0_6_i_ARSIZE <= twiddle_rsc_0_6_ARSIZE;
  twiddle_rsc_0_6_i_ARBURST <= twiddle_rsc_0_6_ARBURST;
  twiddle_rsc_0_6_i_ARCACHE <= twiddle_rsc_0_6_ARCACHE;
  twiddle_rsc_0_6_i_ARPROT <= twiddle_rsc_0_6_ARPROT;
  twiddle_rsc_0_6_i_ARQOS <= twiddle_rsc_0_6_ARQOS;
  twiddle_rsc_0_6_i_ARREGION <= twiddle_rsc_0_6_ARREGION;
  twiddle_rsc_0_6_i_ARUSER(0) <= twiddle_rsc_0_6_ARUSER;
  twiddle_rsc_0_6_RID <= twiddle_rsc_0_6_i_RID(0);
  twiddle_rsc_0_6_RDATA <= twiddle_rsc_0_6_i_RDATA;
  twiddle_rsc_0_6_RRESP <= twiddle_rsc_0_6_i_RRESP;
  twiddle_rsc_0_6_RUSER <= twiddle_rsc_0_6_i_RUSER(0);
  twiddle_rsc_0_6_i_s_raddr_1 <= twiddle_rsc_0_6_i_s_raddr;
  twiddle_rsc_0_6_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_6_i_s_din <= twiddle_rsc_0_6_i_s_din_1;
  twiddle_rsc_0_6_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_6_i_oswt => twiddle_rsc_0_6_i_oswt,
      twiddle_rsc_0_6_i_biwt => twiddle_rsc_0_6_i_biwt,
      twiddle_rsc_0_6_i_bdwt => twiddle_rsc_0_6_i_bdwt,
      twiddle_rsc_0_6_i_bcwt => twiddle_rsc_0_6_i_bcwt,
      twiddle_rsc_0_6_i_s_re_core_sct => twiddle_rsc_0_6_i_s_re_core_sct,
      twiddle_rsc_0_6_i_s_rrdy => twiddle_rsc_0_6_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_6_i_oswt => twiddle_rsc_0_6_i_oswt,
      twiddle_rsc_0_6_i_wen_comp => twiddle_rsc_0_6_i_wen_comp,
      twiddle_rsc_0_6_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_s_raddr_core,
      twiddle_rsc_0_6_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_s_din_mxwt,
      twiddle_rsc_0_6_i_biwt => twiddle_rsc_0_6_i_biwt,
      twiddle_rsc_0_6_i_bdwt => twiddle_rsc_0_6_i_bdwt,
      twiddle_rsc_0_6_i_bcwt => twiddle_rsc_0_6_i_bcwt,
      twiddle_rsc_0_6_i_s_raddr => peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_s_raddr,
      twiddle_rsc_0_6_i_s_raddr_core_sct => twiddle_rsc_0_6_i_s_re_core_sct,
      twiddle_rsc_0_6_i_s_din => peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_6_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_6_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_s_din_mxwt;
  twiddle_rsc_0_6_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_6_i_twiddle_rsc_0_6_wait_dp_inst_twiddle_rsc_0_6_i_s_din
      <= twiddle_rsc_0_6_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_5_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_5_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_5_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_5_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_5_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_5_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_5_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_5_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_5_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_5_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_RID : OUT STD_LOGIC;
    twiddle_rsc_0_5_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_5_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_5_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_5_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_5_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_5_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_5_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_5_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_5_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_5_ARID : IN STD_LOGIC;
    twiddle_rsc_0_5_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_5_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_5_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_5_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_5_BID : OUT STD_LOGIC;
    twiddle_rsc_0_5_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_5_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_5_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_5_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_5_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_5_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_5_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_5_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_5_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_5_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_5_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_5_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_5_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_5_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_5_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_5_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_5_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_5_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_5_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_5_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_5_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_5_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_5_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_5_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_5_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_5_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_5_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_5_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_5_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_5_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_5_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_5_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_5_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_5_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_5_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_5_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_5_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_5_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_5_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_5_i_AWID,
      AWADDR => twiddle_rsc_0_5_i_AWADDR,
      AWLEN => twiddle_rsc_0_5_i_AWLEN,
      AWSIZE => twiddle_rsc_0_5_i_AWSIZE,
      AWBURST => twiddle_rsc_0_5_i_AWBURST,
      AWLOCK => twiddle_rsc_0_5_AWLOCK,
      AWCACHE => twiddle_rsc_0_5_i_AWCACHE,
      AWPROT => twiddle_rsc_0_5_i_AWPROT,
      AWQOS => twiddle_rsc_0_5_i_AWQOS,
      AWREGION => twiddle_rsc_0_5_i_AWREGION,
      AWUSER => twiddle_rsc_0_5_i_AWUSER,
      AWVALID => twiddle_rsc_0_5_AWVALID,
      AWREADY => twiddle_rsc_0_5_AWREADY,
      WDATA => twiddle_rsc_0_5_i_WDATA,
      WSTRB => twiddle_rsc_0_5_i_WSTRB,
      WLAST => twiddle_rsc_0_5_WLAST,
      WUSER => twiddle_rsc_0_5_i_WUSER,
      WVALID => twiddle_rsc_0_5_WVALID,
      WREADY => twiddle_rsc_0_5_WREADY,
      BID => twiddle_rsc_0_5_i_BID,
      BRESP => twiddle_rsc_0_5_i_BRESP,
      BUSER => twiddle_rsc_0_5_i_BUSER,
      BVALID => twiddle_rsc_0_5_BVALID,
      BREADY => twiddle_rsc_0_5_BREADY,
      ARID => twiddle_rsc_0_5_i_ARID,
      ARADDR => twiddle_rsc_0_5_i_ARADDR,
      ARLEN => twiddle_rsc_0_5_i_ARLEN,
      ARSIZE => twiddle_rsc_0_5_i_ARSIZE,
      ARBURST => twiddle_rsc_0_5_i_ARBURST,
      ARLOCK => twiddle_rsc_0_5_ARLOCK,
      ARCACHE => twiddle_rsc_0_5_i_ARCACHE,
      ARPROT => twiddle_rsc_0_5_i_ARPROT,
      ARQOS => twiddle_rsc_0_5_i_ARQOS,
      ARREGION => twiddle_rsc_0_5_i_ARREGION,
      ARUSER => twiddle_rsc_0_5_i_ARUSER,
      ARVALID => twiddle_rsc_0_5_ARVALID,
      ARREADY => twiddle_rsc_0_5_ARREADY,
      RID => twiddle_rsc_0_5_i_RID,
      RDATA => twiddle_rsc_0_5_i_RDATA,
      RRESP => twiddle_rsc_0_5_i_RRESP,
      RLAST => twiddle_rsc_0_5_RLAST,
      RUSER => twiddle_rsc_0_5_i_RUSER,
      RVALID => twiddle_rsc_0_5_RVALID,
      RREADY => twiddle_rsc_0_5_RREADY,
      s_re => twiddle_rsc_0_5_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_5_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_5_i_s_waddr,
      s_din => twiddle_rsc_0_5_i_s_din_1,
      s_dout => twiddle_rsc_0_5_i_s_dout,
      s_rrdy => twiddle_rsc_0_5_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_5_i_s_wrdy,
      is_idle => twiddle_rsc_0_5_is_idle,
      tr_write_done => twiddle_rsc_0_5_tr_write_done,
      s_tdone => twiddle_rsc_0_5_s_tdone
    );
  twiddle_rsc_0_5_i_AWID(0) <= twiddle_rsc_0_5_AWID;
  twiddle_rsc_0_5_i_AWADDR <= twiddle_rsc_0_5_AWADDR;
  twiddle_rsc_0_5_i_AWLEN <= twiddle_rsc_0_5_AWLEN;
  twiddle_rsc_0_5_i_AWSIZE <= twiddle_rsc_0_5_AWSIZE;
  twiddle_rsc_0_5_i_AWBURST <= twiddle_rsc_0_5_AWBURST;
  twiddle_rsc_0_5_i_AWCACHE <= twiddle_rsc_0_5_AWCACHE;
  twiddle_rsc_0_5_i_AWPROT <= twiddle_rsc_0_5_AWPROT;
  twiddle_rsc_0_5_i_AWQOS <= twiddle_rsc_0_5_AWQOS;
  twiddle_rsc_0_5_i_AWREGION <= twiddle_rsc_0_5_AWREGION;
  twiddle_rsc_0_5_i_AWUSER(0) <= twiddle_rsc_0_5_AWUSER;
  twiddle_rsc_0_5_i_WDATA <= twiddle_rsc_0_5_WDATA;
  twiddle_rsc_0_5_i_WSTRB <= twiddle_rsc_0_5_WSTRB;
  twiddle_rsc_0_5_i_WUSER(0) <= twiddle_rsc_0_5_WUSER;
  twiddle_rsc_0_5_BID <= twiddle_rsc_0_5_i_BID(0);
  twiddle_rsc_0_5_BRESP <= twiddle_rsc_0_5_i_BRESP;
  twiddle_rsc_0_5_BUSER <= twiddle_rsc_0_5_i_BUSER(0);
  twiddle_rsc_0_5_i_ARID(0) <= twiddle_rsc_0_5_ARID;
  twiddle_rsc_0_5_i_ARADDR <= twiddle_rsc_0_5_ARADDR;
  twiddle_rsc_0_5_i_ARLEN <= twiddle_rsc_0_5_ARLEN;
  twiddle_rsc_0_5_i_ARSIZE <= twiddle_rsc_0_5_ARSIZE;
  twiddle_rsc_0_5_i_ARBURST <= twiddle_rsc_0_5_ARBURST;
  twiddle_rsc_0_5_i_ARCACHE <= twiddle_rsc_0_5_ARCACHE;
  twiddle_rsc_0_5_i_ARPROT <= twiddle_rsc_0_5_ARPROT;
  twiddle_rsc_0_5_i_ARQOS <= twiddle_rsc_0_5_ARQOS;
  twiddle_rsc_0_5_i_ARREGION <= twiddle_rsc_0_5_ARREGION;
  twiddle_rsc_0_5_i_ARUSER(0) <= twiddle_rsc_0_5_ARUSER;
  twiddle_rsc_0_5_RID <= twiddle_rsc_0_5_i_RID(0);
  twiddle_rsc_0_5_RDATA <= twiddle_rsc_0_5_i_RDATA;
  twiddle_rsc_0_5_RRESP <= twiddle_rsc_0_5_i_RRESP;
  twiddle_rsc_0_5_RUSER <= twiddle_rsc_0_5_i_RUSER(0);
  twiddle_rsc_0_5_i_s_raddr_1 <= twiddle_rsc_0_5_i_s_raddr;
  twiddle_rsc_0_5_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_5_i_s_din <= twiddle_rsc_0_5_i_s_din_1;
  twiddle_rsc_0_5_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_5_i_oswt => twiddle_rsc_0_5_i_oswt,
      twiddle_rsc_0_5_i_biwt => twiddle_rsc_0_5_i_biwt,
      twiddle_rsc_0_5_i_bdwt => twiddle_rsc_0_5_i_bdwt,
      twiddle_rsc_0_5_i_bcwt => twiddle_rsc_0_5_i_bcwt,
      twiddle_rsc_0_5_i_s_re_core_sct => twiddle_rsc_0_5_i_s_re_core_sct,
      twiddle_rsc_0_5_i_s_rrdy => twiddle_rsc_0_5_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_5_i_oswt => twiddle_rsc_0_5_i_oswt,
      twiddle_rsc_0_5_i_wen_comp => twiddle_rsc_0_5_i_wen_comp,
      twiddle_rsc_0_5_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_s_raddr_core,
      twiddle_rsc_0_5_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_s_din_mxwt,
      twiddle_rsc_0_5_i_biwt => twiddle_rsc_0_5_i_biwt,
      twiddle_rsc_0_5_i_bdwt => twiddle_rsc_0_5_i_bdwt,
      twiddle_rsc_0_5_i_bcwt => twiddle_rsc_0_5_i_bcwt,
      twiddle_rsc_0_5_i_s_raddr => peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_s_raddr,
      twiddle_rsc_0_5_i_s_raddr_core_sct => twiddle_rsc_0_5_i_s_re_core_sct,
      twiddle_rsc_0_5_i_s_din => peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_5_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_5_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_s_din_mxwt;
  twiddle_rsc_0_5_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_5_i_twiddle_rsc_0_5_wait_dp_inst_twiddle_rsc_0_5_i_s_din
      <= twiddle_rsc_0_5_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_4_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_4_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_4_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_4_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_4_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_4_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_4_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_4_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_4_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_4_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_RID : OUT STD_LOGIC;
    twiddle_rsc_0_4_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_4_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_4_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_4_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_4_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_4_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_4_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_4_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_4_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_4_ARID : IN STD_LOGIC;
    twiddle_rsc_0_4_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_4_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_4_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_4_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_4_BID : OUT STD_LOGIC;
    twiddle_rsc_0_4_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_4_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_4_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_4_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_4_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_4_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_4_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_4_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_4_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_4_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_4_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_4_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_4_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_4_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_4_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_4_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_4_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_4_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_4_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_4_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_4_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_4_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_4_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_4_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_4_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_4_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_4_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_4_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_4_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_4_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_4_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_4_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_4_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_4_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_4_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_4_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_4_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_4_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_4_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_4_i_AWID,
      AWADDR => twiddle_rsc_0_4_i_AWADDR,
      AWLEN => twiddle_rsc_0_4_i_AWLEN,
      AWSIZE => twiddle_rsc_0_4_i_AWSIZE,
      AWBURST => twiddle_rsc_0_4_i_AWBURST,
      AWLOCK => twiddle_rsc_0_4_AWLOCK,
      AWCACHE => twiddle_rsc_0_4_i_AWCACHE,
      AWPROT => twiddle_rsc_0_4_i_AWPROT,
      AWQOS => twiddle_rsc_0_4_i_AWQOS,
      AWREGION => twiddle_rsc_0_4_i_AWREGION,
      AWUSER => twiddle_rsc_0_4_i_AWUSER,
      AWVALID => twiddle_rsc_0_4_AWVALID,
      AWREADY => twiddle_rsc_0_4_AWREADY,
      WDATA => twiddle_rsc_0_4_i_WDATA,
      WSTRB => twiddle_rsc_0_4_i_WSTRB,
      WLAST => twiddle_rsc_0_4_WLAST,
      WUSER => twiddle_rsc_0_4_i_WUSER,
      WVALID => twiddle_rsc_0_4_WVALID,
      WREADY => twiddle_rsc_0_4_WREADY,
      BID => twiddle_rsc_0_4_i_BID,
      BRESP => twiddle_rsc_0_4_i_BRESP,
      BUSER => twiddle_rsc_0_4_i_BUSER,
      BVALID => twiddle_rsc_0_4_BVALID,
      BREADY => twiddle_rsc_0_4_BREADY,
      ARID => twiddle_rsc_0_4_i_ARID,
      ARADDR => twiddle_rsc_0_4_i_ARADDR,
      ARLEN => twiddle_rsc_0_4_i_ARLEN,
      ARSIZE => twiddle_rsc_0_4_i_ARSIZE,
      ARBURST => twiddle_rsc_0_4_i_ARBURST,
      ARLOCK => twiddle_rsc_0_4_ARLOCK,
      ARCACHE => twiddle_rsc_0_4_i_ARCACHE,
      ARPROT => twiddle_rsc_0_4_i_ARPROT,
      ARQOS => twiddle_rsc_0_4_i_ARQOS,
      ARREGION => twiddle_rsc_0_4_i_ARREGION,
      ARUSER => twiddle_rsc_0_4_i_ARUSER,
      ARVALID => twiddle_rsc_0_4_ARVALID,
      ARREADY => twiddle_rsc_0_4_ARREADY,
      RID => twiddle_rsc_0_4_i_RID,
      RDATA => twiddle_rsc_0_4_i_RDATA,
      RRESP => twiddle_rsc_0_4_i_RRESP,
      RLAST => twiddle_rsc_0_4_RLAST,
      RUSER => twiddle_rsc_0_4_i_RUSER,
      RVALID => twiddle_rsc_0_4_RVALID,
      RREADY => twiddle_rsc_0_4_RREADY,
      s_re => twiddle_rsc_0_4_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_4_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_4_i_s_waddr,
      s_din => twiddle_rsc_0_4_i_s_din_1,
      s_dout => twiddle_rsc_0_4_i_s_dout,
      s_rrdy => twiddle_rsc_0_4_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_4_i_s_wrdy,
      is_idle => twiddle_rsc_0_4_is_idle,
      tr_write_done => twiddle_rsc_0_4_tr_write_done,
      s_tdone => twiddle_rsc_0_4_s_tdone
    );
  twiddle_rsc_0_4_i_AWID(0) <= twiddle_rsc_0_4_AWID;
  twiddle_rsc_0_4_i_AWADDR <= twiddle_rsc_0_4_AWADDR;
  twiddle_rsc_0_4_i_AWLEN <= twiddle_rsc_0_4_AWLEN;
  twiddle_rsc_0_4_i_AWSIZE <= twiddle_rsc_0_4_AWSIZE;
  twiddle_rsc_0_4_i_AWBURST <= twiddle_rsc_0_4_AWBURST;
  twiddle_rsc_0_4_i_AWCACHE <= twiddle_rsc_0_4_AWCACHE;
  twiddle_rsc_0_4_i_AWPROT <= twiddle_rsc_0_4_AWPROT;
  twiddle_rsc_0_4_i_AWQOS <= twiddle_rsc_0_4_AWQOS;
  twiddle_rsc_0_4_i_AWREGION <= twiddle_rsc_0_4_AWREGION;
  twiddle_rsc_0_4_i_AWUSER(0) <= twiddle_rsc_0_4_AWUSER;
  twiddle_rsc_0_4_i_WDATA <= twiddle_rsc_0_4_WDATA;
  twiddle_rsc_0_4_i_WSTRB <= twiddle_rsc_0_4_WSTRB;
  twiddle_rsc_0_4_i_WUSER(0) <= twiddle_rsc_0_4_WUSER;
  twiddle_rsc_0_4_BID <= twiddle_rsc_0_4_i_BID(0);
  twiddle_rsc_0_4_BRESP <= twiddle_rsc_0_4_i_BRESP;
  twiddle_rsc_0_4_BUSER <= twiddle_rsc_0_4_i_BUSER(0);
  twiddle_rsc_0_4_i_ARID(0) <= twiddle_rsc_0_4_ARID;
  twiddle_rsc_0_4_i_ARADDR <= twiddle_rsc_0_4_ARADDR;
  twiddle_rsc_0_4_i_ARLEN <= twiddle_rsc_0_4_ARLEN;
  twiddle_rsc_0_4_i_ARSIZE <= twiddle_rsc_0_4_ARSIZE;
  twiddle_rsc_0_4_i_ARBURST <= twiddle_rsc_0_4_ARBURST;
  twiddle_rsc_0_4_i_ARCACHE <= twiddle_rsc_0_4_ARCACHE;
  twiddle_rsc_0_4_i_ARPROT <= twiddle_rsc_0_4_ARPROT;
  twiddle_rsc_0_4_i_ARQOS <= twiddle_rsc_0_4_ARQOS;
  twiddle_rsc_0_4_i_ARREGION <= twiddle_rsc_0_4_ARREGION;
  twiddle_rsc_0_4_i_ARUSER(0) <= twiddle_rsc_0_4_ARUSER;
  twiddle_rsc_0_4_RID <= twiddle_rsc_0_4_i_RID(0);
  twiddle_rsc_0_4_RDATA <= twiddle_rsc_0_4_i_RDATA;
  twiddle_rsc_0_4_RRESP <= twiddle_rsc_0_4_i_RRESP;
  twiddle_rsc_0_4_RUSER <= twiddle_rsc_0_4_i_RUSER(0);
  twiddle_rsc_0_4_i_s_raddr_1 <= twiddle_rsc_0_4_i_s_raddr;
  twiddle_rsc_0_4_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_4_i_s_din <= twiddle_rsc_0_4_i_s_din_1;
  twiddle_rsc_0_4_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_4_i_oswt => twiddle_rsc_0_4_i_oswt,
      twiddle_rsc_0_4_i_biwt => twiddle_rsc_0_4_i_biwt,
      twiddle_rsc_0_4_i_bdwt => twiddle_rsc_0_4_i_bdwt,
      twiddle_rsc_0_4_i_bcwt => twiddle_rsc_0_4_i_bcwt,
      twiddle_rsc_0_4_i_s_re_core_sct => twiddle_rsc_0_4_i_s_re_core_sct,
      twiddle_rsc_0_4_i_s_rrdy => twiddle_rsc_0_4_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_4_i_oswt => twiddle_rsc_0_4_i_oswt,
      twiddle_rsc_0_4_i_wen_comp => twiddle_rsc_0_4_i_wen_comp,
      twiddle_rsc_0_4_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_s_raddr_core,
      twiddle_rsc_0_4_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_s_din_mxwt,
      twiddle_rsc_0_4_i_biwt => twiddle_rsc_0_4_i_biwt,
      twiddle_rsc_0_4_i_bdwt => twiddle_rsc_0_4_i_bdwt,
      twiddle_rsc_0_4_i_bcwt => twiddle_rsc_0_4_i_bcwt,
      twiddle_rsc_0_4_i_s_raddr => peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_s_raddr,
      twiddle_rsc_0_4_i_s_raddr_core_sct => twiddle_rsc_0_4_i_s_re_core_sct,
      twiddle_rsc_0_4_i_s_din => peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_4_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_4_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_s_din_mxwt;
  twiddle_rsc_0_4_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_4_i_twiddle_rsc_0_4_wait_dp_inst_twiddle_rsc_0_4_i_s_din
      <= twiddle_rsc_0_4_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_3_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_3_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_3_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_3_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_3_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_3_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_3_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_3_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_3_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_3_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_RID : OUT STD_LOGIC;
    twiddle_rsc_0_3_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_3_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_3_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_3_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_3_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_3_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_3_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_3_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_3_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_3_ARID : IN STD_LOGIC;
    twiddle_rsc_0_3_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_3_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_3_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_3_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_3_BID : OUT STD_LOGIC;
    twiddle_rsc_0_3_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_3_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_3_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_3_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_3_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_3_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_3_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_3_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_3_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_3_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_3_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_3_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_3_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_3_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_3_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_3_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_3_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_3_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_3_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_3_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_3_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_3_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_3_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_3_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_3_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_3_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_3_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_3_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_3_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_3_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_3_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_3_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_3_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_3_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_3_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_3_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_3_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_3_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_3_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_3_i_AWID,
      AWADDR => twiddle_rsc_0_3_i_AWADDR,
      AWLEN => twiddle_rsc_0_3_i_AWLEN,
      AWSIZE => twiddle_rsc_0_3_i_AWSIZE,
      AWBURST => twiddle_rsc_0_3_i_AWBURST,
      AWLOCK => twiddle_rsc_0_3_AWLOCK,
      AWCACHE => twiddle_rsc_0_3_i_AWCACHE,
      AWPROT => twiddle_rsc_0_3_i_AWPROT,
      AWQOS => twiddle_rsc_0_3_i_AWQOS,
      AWREGION => twiddle_rsc_0_3_i_AWREGION,
      AWUSER => twiddle_rsc_0_3_i_AWUSER,
      AWVALID => twiddle_rsc_0_3_AWVALID,
      AWREADY => twiddle_rsc_0_3_AWREADY,
      WDATA => twiddle_rsc_0_3_i_WDATA,
      WSTRB => twiddle_rsc_0_3_i_WSTRB,
      WLAST => twiddle_rsc_0_3_WLAST,
      WUSER => twiddle_rsc_0_3_i_WUSER,
      WVALID => twiddle_rsc_0_3_WVALID,
      WREADY => twiddle_rsc_0_3_WREADY,
      BID => twiddle_rsc_0_3_i_BID,
      BRESP => twiddle_rsc_0_3_i_BRESP,
      BUSER => twiddle_rsc_0_3_i_BUSER,
      BVALID => twiddle_rsc_0_3_BVALID,
      BREADY => twiddle_rsc_0_3_BREADY,
      ARID => twiddle_rsc_0_3_i_ARID,
      ARADDR => twiddle_rsc_0_3_i_ARADDR,
      ARLEN => twiddle_rsc_0_3_i_ARLEN,
      ARSIZE => twiddle_rsc_0_3_i_ARSIZE,
      ARBURST => twiddle_rsc_0_3_i_ARBURST,
      ARLOCK => twiddle_rsc_0_3_ARLOCK,
      ARCACHE => twiddle_rsc_0_3_i_ARCACHE,
      ARPROT => twiddle_rsc_0_3_i_ARPROT,
      ARQOS => twiddle_rsc_0_3_i_ARQOS,
      ARREGION => twiddle_rsc_0_3_i_ARREGION,
      ARUSER => twiddle_rsc_0_3_i_ARUSER,
      ARVALID => twiddle_rsc_0_3_ARVALID,
      ARREADY => twiddle_rsc_0_3_ARREADY,
      RID => twiddle_rsc_0_3_i_RID,
      RDATA => twiddle_rsc_0_3_i_RDATA,
      RRESP => twiddle_rsc_0_3_i_RRESP,
      RLAST => twiddle_rsc_0_3_RLAST,
      RUSER => twiddle_rsc_0_3_i_RUSER,
      RVALID => twiddle_rsc_0_3_RVALID,
      RREADY => twiddle_rsc_0_3_RREADY,
      s_re => twiddle_rsc_0_3_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_3_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_3_i_s_waddr,
      s_din => twiddle_rsc_0_3_i_s_din_1,
      s_dout => twiddle_rsc_0_3_i_s_dout,
      s_rrdy => twiddle_rsc_0_3_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_3_i_s_wrdy,
      is_idle => twiddle_rsc_0_3_is_idle,
      tr_write_done => twiddle_rsc_0_3_tr_write_done,
      s_tdone => twiddle_rsc_0_3_s_tdone
    );
  twiddle_rsc_0_3_i_AWID(0) <= twiddle_rsc_0_3_AWID;
  twiddle_rsc_0_3_i_AWADDR <= twiddle_rsc_0_3_AWADDR;
  twiddle_rsc_0_3_i_AWLEN <= twiddle_rsc_0_3_AWLEN;
  twiddle_rsc_0_3_i_AWSIZE <= twiddle_rsc_0_3_AWSIZE;
  twiddle_rsc_0_3_i_AWBURST <= twiddle_rsc_0_3_AWBURST;
  twiddle_rsc_0_3_i_AWCACHE <= twiddle_rsc_0_3_AWCACHE;
  twiddle_rsc_0_3_i_AWPROT <= twiddle_rsc_0_3_AWPROT;
  twiddle_rsc_0_3_i_AWQOS <= twiddle_rsc_0_3_AWQOS;
  twiddle_rsc_0_3_i_AWREGION <= twiddle_rsc_0_3_AWREGION;
  twiddle_rsc_0_3_i_AWUSER(0) <= twiddle_rsc_0_3_AWUSER;
  twiddle_rsc_0_3_i_WDATA <= twiddle_rsc_0_3_WDATA;
  twiddle_rsc_0_3_i_WSTRB <= twiddle_rsc_0_3_WSTRB;
  twiddle_rsc_0_3_i_WUSER(0) <= twiddle_rsc_0_3_WUSER;
  twiddle_rsc_0_3_BID <= twiddle_rsc_0_3_i_BID(0);
  twiddle_rsc_0_3_BRESP <= twiddle_rsc_0_3_i_BRESP;
  twiddle_rsc_0_3_BUSER <= twiddle_rsc_0_3_i_BUSER(0);
  twiddle_rsc_0_3_i_ARID(0) <= twiddle_rsc_0_3_ARID;
  twiddle_rsc_0_3_i_ARADDR <= twiddle_rsc_0_3_ARADDR;
  twiddle_rsc_0_3_i_ARLEN <= twiddle_rsc_0_3_ARLEN;
  twiddle_rsc_0_3_i_ARSIZE <= twiddle_rsc_0_3_ARSIZE;
  twiddle_rsc_0_3_i_ARBURST <= twiddle_rsc_0_3_ARBURST;
  twiddle_rsc_0_3_i_ARCACHE <= twiddle_rsc_0_3_ARCACHE;
  twiddle_rsc_0_3_i_ARPROT <= twiddle_rsc_0_3_ARPROT;
  twiddle_rsc_0_3_i_ARQOS <= twiddle_rsc_0_3_ARQOS;
  twiddle_rsc_0_3_i_ARREGION <= twiddle_rsc_0_3_ARREGION;
  twiddle_rsc_0_3_i_ARUSER(0) <= twiddle_rsc_0_3_ARUSER;
  twiddle_rsc_0_3_RID <= twiddle_rsc_0_3_i_RID(0);
  twiddle_rsc_0_3_RDATA <= twiddle_rsc_0_3_i_RDATA;
  twiddle_rsc_0_3_RRESP <= twiddle_rsc_0_3_i_RRESP;
  twiddle_rsc_0_3_RUSER <= twiddle_rsc_0_3_i_RUSER(0);
  twiddle_rsc_0_3_i_s_raddr_1 <= twiddle_rsc_0_3_i_s_raddr;
  twiddle_rsc_0_3_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_3_i_s_din <= twiddle_rsc_0_3_i_s_din_1;
  twiddle_rsc_0_3_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_3_i_oswt => twiddle_rsc_0_3_i_oswt,
      twiddle_rsc_0_3_i_biwt => twiddle_rsc_0_3_i_biwt,
      twiddle_rsc_0_3_i_bdwt => twiddle_rsc_0_3_i_bdwt,
      twiddle_rsc_0_3_i_bcwt => twiddle_rsc_0_3_i_bcwt,
      twiddle_rsc_0_3_i_s_re_core_sct => twiddle_rsc_0_3_i_s_re_core_sct,
      twiddle_rsc_0_3_i_s_rrdy => twiddle_rsc_0_3_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_3_i_oswt => twiddle_rsc_0_3_i_oswt,
      twiddle_rsc_0_3_i_wen_comp => twiddle_rsc_0_3_i_wen_comp,
      twiddle_rsc_0_3_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_s_raddr_core,
      twiddle_rsc_0_3_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_s_din_mxwt,
      twiddle_rsc_0_3_i_biwt => twiddle_rsc_0_3_i_biwt,
      twiddle_rsc_0_3_i_bdwt => twiddle_rsc_0_3_i_bdwt,
      twiddle_rsc_0_3_i_bcwt => twiddle_rsc_0_3_i_bcwt,
      twiddle_rsc_0_3_i_s_raddr => peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_s_raddr,
      twiddle_rsc_0_3_i_s_raddr_core_sct => twiddle_rsc_0_3_i_s_re_core_sct,
      twiddle_rsc_0_3_i_s_din => peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_3_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_3_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_s_din_mxwt;
  twiddle_rsc_0_3_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_3_i_twiddle_rsc_0_3_wait_dp_inst_twiddle_rsc_0_3_i_s_din
      <= twiddle_rsc_0_3_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_2_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_2_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_2_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_2_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_2_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_2_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_2_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_2_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_2_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_2_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_RID : OUT STD_LOGIC;
    twiddle_rsc_0_2_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_2_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_2_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_2_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_2_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_2_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_2_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_2_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_2_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_2_ARID : IN STD_LOGIC;
    twiddle_rsc_0_2_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_2_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_2_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_2_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_2_BID : OUT STD_LOGIC;
    twiddle_rsc_0_2_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_2_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_2_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_2_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_2_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_2_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_2_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_2_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_2_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_2_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_2_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_2_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_2_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_2_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_2_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_2_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_2_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_2_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_2_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_2_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_2_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_2_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_2_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_2_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_2_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_2_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_2_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_2_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_2_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_2_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_2_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_2_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_2_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_2_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_2_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_2_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_2_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_2_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_2_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_2_i_AWID,
      AWADDR => twiddle_rsc_0_2_i_AWADDR,
      AWLEN => twiddle_rsc_0_2_i_AWLEN,
      AWSIZE => twiddle_rsc_0_2_i_AWSIZE,
      AWBURST => twiddle_rsc_0_2_i_AWBURST,
      AWLOCK => twiddle_rsc_0_2_AWLOCK,
      AWCACHE => twiddle_rsc_0_2_i_AWCACHE,
      AWPROT => twiddle_rsc_0_2_i_AWPROT,
      AWQOS => twiddle_rsc_0_2_i_AWQOS,
      AWREGION => twiddle_rsc_0_2_i_AWREGION,
      AWUSER => twiddle_rsc_0_2_i_AWUSER,
      AWVALID => twiddle_rsc_0_2_AWVALID,
      AWREADY => twiddle_rsc_0_2_AWREADY,
      WDATA => twiddle_rsc_0_2_i_WDATA,
      WSTRB => twiddle_rsc_0_2_i_WSTRB,
      WLAST => twiddle_rsc_0_2_WLAST,
      WUSER => twiddle_rsc_0_2_i_WUSER,
      WVALID => twiddle_rsc_0_2_WVALID,
      WREADY => twiddle_rsc_0_2_WREADY,
      BID => twiddle_rsc_0_2_i_BID,
      BRESP => twiddle_rsc_0_2_i_BRESP,
      BUSER => twiddle_rsc_0_2_i_BUSER,
      BVALID => twiddle_rsc_0_2_BVALID,
      BREADY => twiddle_rsc_0_2_BREADY,
      ARID => twiddle_rsc_0_2_i_ARID,
      ARADDR => twiddle_rsc_0_2_i_ARADDR,
      ARLEN => twiddle_rsc_0_2_i_ARLEN,
      ARSIZE => twiddle_rsc_0_2_i_ARSIZE,
      ARBURST => twiddle_rsc_0_2_i_ARBURST,
      ARLOCK => twiddle_rsc_0_2_ARLOCK,
      ARCACHE => twiddle_rsc_0_2_i_ARCACHE,
      ARPROT => twiddle_rsc_0_2_i_ARPROT,
      ARQOS => twiddle_rsc_0_2_i_ARQOS,
      ARREGION => twiddle_rsc_0_2_i_ARREGION,
      ARUSER => twiddle_rsc_0_2_i_ARUSER,
      ARVALID => twiddle_rsc_0_2_ARVALID,
      ARREADY => twiddle_rsc_0_2_ARREADY,
      RID => twiddle_rsc_0_2_i_RID,
      RDATA => twiddle_rsc_0_2_i_RDATA,
      RRESP => twiddle_rsc_0_2_i_RRESP,
      RLAST => twiddle_rsc_0_2_RLAST,
      RUSER => twiddle_rsc_0_2_i_RUSER,
      RVALID => twiddle_rsc_0_2_RVALID,
      RREADY => twiddle_rsc_0_2_RREADY,
      s_re => twiddle_rsc_0_2_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_2_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_2_i_s_waddr,
      s_din => twiddle_rsc_0_2_i_s_din_1,
      s_dout => twiddle_rsc_0_2_i_s_dout,
      s_rrdy => twiddle_rsc_0_2_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_2_i_s_wrdy,
      is_idle => twiddle_rsc_0_2_is_idle,
      tr_write_done => twiddle_rsc_0_2_tr_write_done,
      s_tdone => twiddle_rsc_0_2_s_tdone
    );
  twiddle_rsc_0_2_i_AWID(0) <= twiddle_rsc_0_2_AWID;
  twiddle_rsc_0_2_i_AWADDR <= twiddle_rsc_0_2_AWADDR;
  twiddle_rsc_0_2_i_AWLEN <= twiddle_rsc_0_2_AWLEN;
  twiddle_rsc_0_2_i_AWSIZE <= twiddle_rsc_0_2_AWSIZE;
  twiddle_rsc_0_2_i_AWBURST <= twiddle_rsc_0_2_AWBURST;
  twiddle_rsc_0_2_i_AWCACHE <= twiddle_rsc_0_2_AWCACHE;
  twiddle_rsc_0_2_i_AWPROT <= twiddle_rsc_0_2_AWPROT;
  twiddle_rsc_0_2_i_AWQOS <= twiddle_rsc_0_2_AWQOS;
  twiddle_rsc_0_2_i_AWREGION <= twiddle_rsc_0_2_AWREGION;
  twiddle_rsc_0_2_i_AWUSER(0) <= twiddle_rsc_0_2_AWUSER;
  twiddle_rsc_0_2_i_WDATA <= twiddle_rsc_0_2_WDATA;
  twiddle_rsc_0_2_i_WSTRB <= twiddle_rsc_0_2_WSTRB;
  twiddle_rsc_0_2_i_WUSER(0) <= twiddle_rsc_0_2_WUSER;
  twiddle_rsc_0_2_BID <= twiddle_rsc_0_2_i_BID(0);
  twiddle_rsc_0_2_BRESP <= twiddle_rsc_0_2_i_BRESP;
  twiddle_rsc_0_2_BUSER <= twiddle_rsc_0_2_i_BUSER(0);
  twiddle_rsc_0_2_i_ARID(0) <= twiddle_rsc_0_2_ARID;
  twiddle_rsc_0_2_i_ARADDR <= twiddle_rsc_0_2_ARADDR;
  twiddle_rsc_0_2_i_ARLEN <= twiddle_rsc_0_2_ARLEN;
  twiddle_rsc_0_2_i_ARSIZE <= twiddle_rsc_0_2_ARSIZE;
  twiddle_rsc_0_2_i_ARBURST <= twiddle_rsc_0_2_ARBURST;
  twiddle_rsc_0_2_i_ARCACHE <= twiddle_rsc_0_2_ARCACHE;
  twiddle_rsc_0_2_i_ARPROT <= twiddle_rsc_0_2_ARPROT;
  twiddle_rsc_0_2_i_ARQOS <= twiddle_rsc_0_2_ARQOS;
  twiddle_rsc_0_2_i_ARREGION <= twiddle_rsc_0_2_ARREGION;
  twiddle_rsc_0_2_i_ARUSER(0) <= twiddle_rsc_0_2_ARUSER;
  twiddle_rsc_0_2_RID <= twiddle_rsc_0_2_i_RID(0);
  twiddle_rsc_0_2_RDATA <= twiddle_rsc_0_2_i_RDATA;
  twiddle_rsc_0_2_RRESP <= twiddle_rsc_0_2_i_RRESP;
  twiddle_rsc_0_2_RUSER <= twiddle_rsc_0_2_i_RUSER(0);
  twiddle_rsc_0_2_i_s_raddr_1 <= twiddle_rsc_0_2_i_s_raddr;
  twiddle_rsc_0_2_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_2_i_s_din <= twiddle_rsc_0_2_i_s_din_1;
  twiddle_rsc_0_2_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_2_i_oswt => twiddle_rsc_0_2_i_oswt,
      twiddle_rsc_0_2_i_biwt => twiddle_rsc_0_2_i_biwt,
      twiddle_rsc_0_2_i_bdwt => twiddle_rsc_0_2_i_bdwt,
      twiddle_rsc_0_2_i_bcwt => twiddle_rsc_0_2_i_bcwt,
      twiddle_rsc_0_2_i_s_re_core_sct => twiddle_rsc_0_2_i_s_re_core_sct,
      twiddle_rsc_0_2_i_s_rrdy => twiddle_rsc_0_2_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_2_i_oswt => twiddle_rsc_0_2_i_oswt,
      twiddle_rsc_0_2_i_wen_comp => twiddle_rsc_0_2_i_wen_comp,
      twiddle_rsc_0_2_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_s_raddr_core,
      twiddle_rsc_0_2_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_s_din_mxwt,
      twiddle_rsc_0_2_i_biwt => twiddle_rsc_0_2_i_biwt,
      twiddle_rsc_0_2_i_bdwt => twiddle_rsc_0_2_i_bdwt,
      twiddle_rsc_0_2_i_bcwt => twiddle_rsc_0_2_i_bcwt,
      twiddle_rsc_0_2_i_s_raddr => peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_s_raddr,
      twiddle_rsc_0_2_i_s_raddr_core_sct => twiddle_rsc_0_2_i_s_re_core_sct,
      twiddle_rsc_0_2_i_s_din => peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_2_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_2_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_s_din_mxwt;
  twiddle_rsc_0_2_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_2_i_twiddle_rsc_0_2_wait_dp_inst_twiddle_rsc_0_2_i_s_din
      <= twiddle_rsc_0_2_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_1_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_1_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_1_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_1_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_1_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_1_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_1_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_1_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_1_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_1_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_RID : OUT STD_LOGIC;
    twiddle_rsc_0_1_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_1_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_1_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_1_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_1_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_1_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_1_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_1_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_1_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_1_ARID : IN STD_LOGIC;
    twiddle_rsc_0_1_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_1_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_1_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_1_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_1_BID : OUT STD_LOGIC;
    twiddle_rsc_0_1_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_1_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_1_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_1_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_1_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_1_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_1_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_1_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_1_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_1_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_1_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_1_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_1_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_1_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_1_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_1_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_1_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_1_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_1_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_1_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_1_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_1_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_1_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_1_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_1_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_1_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_1_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_1_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_1_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_1_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_1_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_1_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_1_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_1_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_1_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_1_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_1_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_1_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_1_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_1_i_AWID,
      AWADDR => twiddle_rsc_0_1_i_AWADDR,
      AWLEN => twiddle_rsc_0_1_i_AWLEN,
      AWSIZE => twiddle_rsc_0_1_i_AWSIZE,
      AWBURST => twiddle_rsc_0_1_i_AWBURST,
      AWLOCK => twiddle_rsc_0_1_AWLOCK,
      AWCACHE => twiddle_rsc_0_1_i_AWCACHE,
      AWPROT => twiddle_rsc_0_1_i_AWPROT,
      AWQOS => twiddle_rsc_0_1_i_AWQOS,
      AWREGION => twiddle_rsc_0_1_i_AWREGION,
      AWUSER => twiddle_rsc_0_1_i_AWUSER,
      AWVALID => twiddle_rsc_0_1_AWVALID,
      AWREADY => twiddle_rsc_0_1_AWREADY,
      WDATA => twiddle_rsc_0_1_i_WDATA,
      WSTRB => twiddle_rsc_0_1_i_WSTRB,
      WLAST => twiddle_rsc_0_1_WLAST,
      WUSER => twiddle_rsc_0_1_i_WUSER,
      WVALID => twiddle_rsc_0_1_WVALID,
      WREADY => twiddle_rsc_0_1_WREADY,
      BID => twiddle_rsc_0_1_i_BID,
      BRESP => twiddle_rsc_0_1_i_BRESP,
      BUSER => twiddle_rsc_0_1_i_BUSER,
      BVALID => twiddle_rsc_0_1_BVALID,
      BREADY => twiddle_rsc_0_1_BREADY,
      ARID => twiddle_rsc_0_1_i_ARID,
      ARADDR => twiddle_rsc_0_1_i_ARADDR,
      ARLEN => twiddle_rsc_0_1_i_ARLEN,
      ARSIZE => twiddle_rsc_0_1_i_ARSIZE,
      ARBURST => twiddle_rsc_0_1_i_ARBURST,
      ARLOCK => twiddle_rsc_0_1_ARLOCK,
      ARCACHE => twiddle_rsc_0_1_i_ARCACHE,
      ARPROT => twiddle_rsc_0_1_i_ARPROT,
      ARQOS => twiddle_rsc_0_1_i_ARQOS,
      ARREGION => twiddle_rsc_0_1_i_ARREGION,
      ARUSER => twiddle_rsc_0_1_i_ARUSER,
      ARVALID => twiddle_rsc_0_1_ARVALID,
      ARREADY => twiddle_rsc_0_1_ARREADY,
      RID => twiddle_rsc_0_1_i_RID,
      RDATA => twiddle_rsc_0_1_i_RDATA,
      RRESP => twiddle_rsc_0_1_i_RRESP,
      RLAST => twiddle_rsc_0_1_RLAST,
      RUSER => twiddle_rsc_0_1_i_RUSER,
      RVALID => twiddle_rsc_0_1_RVALID,
      RREADY => twiddle_rsc_0_1_RREADY,
      s_re => twiddle_rsc_0_1_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_1_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_1_i_s_waddr,
      s_din => twiddle_rsc_0_1_i_s_din_1,
      s_dout => twiddle_rsc_0_1_i_s_dout,
      s_rrdy => twiddle_rsc_0_1_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_1_i_s_wrdy,
      is_idle => twiddle_rsc_0_1_is_idle,
      tr_write_done => twiddle_rsc_0_1_tr_write_done,
      s_tdone => twiddle_rsc_0_1_s_tdone
    );
  twiddle_rsc_0_1_i_AWID(0) <= twiddle_rsc_0_1_AWID;
  twiddle_rsc_0_1_i_AWADDR <= twiddle_rsc_0_1_AWADDR;
  twiddle_rsc_0_1_i_AWLEN <= twiddle_rsc_0_1_AWLEN;
  twiddle_rsc_0_1_i_AWSIZE <= twiddle_rsc_0_1_AWSIZE;
  twiddle_rsc_0_1_i_AWBURST <= twiddle_rsc_0_1_AWBURST;
  twiddle_rsc_0_1_i_AWCACHE <= twiddle_rsc_0_1_AWCACHE;
  twiddle_rsc_0_1_i_AWPROT <= twiddle_rsc_0_1_AWPROT;
  twiddle_rsc_0_1_i_AWQOS <= twiddle_rsc_0_1_AWQOS;
  twiddle_rsc_0_1_i_AWREGION <= twiddle_rsc_0_1_AWREGION;
  twiddle_rsc_0_1_i_AWUSER(0) <= twiddle_rsc_0_1_AWUSER;
  twiddle_rsc_0_1_i_WDATA <= twiddle_rsc_0_1_WDATA;
  twiddle_rsc_0_1_i_WSTRB <= twiddle_rsc_0_1_WSTRB;
  twiddle_rsc_0_1_i_WUSER(0) <= twiddle_rsc_0_1_WUSER;
  twiddle_rsc_0_1_BID <= twiddle_rsc_0_1_i_BID(0);
  twiddle_rsc_0_1_BRESP <= twiddle_rsc_0_1_i_BRESP;
  twiddle_rsc_0_1_BUSER <= twiddle_rsc_0_1_i_BUSER(0);
  twiddle_rsc_0_1_i_ARID(0) <= twiddle_rsc_0_1_ARID;
  twiddle_rsc_0_1_i_ARADDR <= twiddle_rsc_0_1_ARADDR;
  twiddle_rsc_0_1_i_ARLEN <= twiddle_rsc_0_1_ARLEN;
  twiddle_rsc_0_1_i_ARSIZE <= twiddle_rsc_0_1_ARSIZE;
  twiddle_rsc_0_1_i_ARBURST <= twiddle_rsc_0_1_ARBURST;
  twiddle_rsc_0_1_i_ARCACHE <= twiddle_rsc_0_1_ARCACHE;
  twiddle_rsc_0_1_i_ARPROT <= twiddle_rsc_0_1_ARPROT;
  twiddle_rsc_0_1_i_ARQOS <= twiddle_rsc_0_1_ARQOS;
  twiddle_rsc_0_1_i_ARREGION <= twiddle_rsc_0_1_ARREGION;
  twiddle_rsc_0_1_i_ARUSER(0) <= twiddle_rsc_0_1_ARUSER;
  twiddle_rsc_0_1_RID <= twiddle_rsc_0_1_i_RID(0);
  twiddle_rsc_0_1_RDATA <= twiddle_rsc_0_1_i_RDATA;
  twiddle_rsc_0_1_RRESP <= twiddle_rsc_0_1_i_RRESP;
  twiddle_rsc_0_1_RUSER <= twiddle_rsc_0_1_i_RUSER(0);
  twiddle_rsc_0_1_i_s_raddr_1 <= twiddle_rsc_0_1_i_s_raddr;
  twiddle_rsc_0_1_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_1_i_s_din <= twiddle_rsc_0_1_i_s_din_1;
  twiddle_rsc_0_1_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_1_i_oswt => twiddle_rsc_0_1_i_oswt,
      twiddle_rsc_0_1_i_biwt => twiddle_rsc_0_1_i_biwt,
      twiddle_rsc_0_1_i_bdwt => twiddle_rsc_0_1_i_bdwt,
      twiddle_rsc_0_1_i_bcwt => twiddle_rsc_0_1_i_bcwt,
      twiddle_rsc_0_1_i_s_re_core_sct => twiddle_rsc_0_1_i_s_re_core_sct,
      twiddle_rsc_0_1_i_s_rrdy => twiddle_rsc_0_1_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_1_i_oswt => twiddle_rsc_0_1_i_oswt,
      twiddle_rsc_0_1_i_wen_comp => twiddle_rsc_0_1_i_wen_comp,
      twiddle_rsc_0_1_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_s_raddr_core,
      twiddle_rsc_0_1_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_s_din_mxwt,
      twiddle_rsc_0_1_i_biwt => twiddle_rsc_0_1_i_biwt,
      twiddle_rsc_0_1_i_bdwt => twiddle_rsc_0_1_i_bdwt,
      twiddle_rsc_0_1_i_bcwt => twiddle_rsc_0_1_i_bcwt,
      twiddle_rsc_0_1_i_s_raddr => peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_s_raddr,
      twiddle_rsc_0_1_i_s_raddr_core_sct => twiddle_rsc_0_1_i_s_re_core_sct,
      twiddle_rsc_0_1_i_s_din => peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_1_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_1_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_s_din_mxwt;
  twiddle_rsc_0_1_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_1_i_twiddle_rsc_0_1_wait_dp_inst_twiddle_rsc_0_1_i_s_din
      <= twiddle_rsc_0_1_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_twiddle_rsc_0_0_i
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_twiddle_rsc_0_0_i IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    twiddle_rsc_0_0_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_0_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_0_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_0_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_0_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_0_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_RID : OUT STD_LOGIC;
    twiddle_rsc_0_0_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_0_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_0_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_0_ARID : IN STD_LOGIC;
    twiddle_rsc_0_0_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_0_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_0_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_0_BID : OUT STD_LOGIC;
    twiddle_rsc_0_0_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_0_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_0_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_0_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_0_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_0_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_0_AWID : IN STD_LOGIC;
    core_wen : IN STD_LOGIC;
    twiddle_rsc_0_0_i_oswt : IN STD_LOGIC;
    twiddle_rsc_0_0_i_wen_comp : OUT STD_LOGIC;
    twiddle_rsc_0_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
    twiddle_rsc_0_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
  );
END peaseNTT_core_twiddle_rsc_0_0_i;

ARCHITECTURE v29 OF peaseNTT_core_twiddle_rsc_0_0_i IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL twiddle_rsc_0_0_i_biwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_bdwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_bcwt : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_s_re_core_sct : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_s_raddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_s_din : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_s_rrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_s_wrdy : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_is_idle : STD_LOGIC;

  SIGNAL twiddle_rsc_0_0_i_AWID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_AWUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_WUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_BID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_BUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_ARID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_ARUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_RID : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_RUSER : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_s_raddr_1 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_s_waddr : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_s_din_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_s_dout : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_0_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_0_i_biwt : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_bdwt : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_bcwt : IN STD_LOGIC;
      twiddle_rsc_0_0_i_s_re_core_sct : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_s_rrdy : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_0_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_0_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_0_i_biwt : IN STD_LOGIC;
      twiddle_rsc_0_0_i_bdwt : IN STD_LOGIC;
      twiddle_rsc_0_0_i_bcwt : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_s_raddr : OUT STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_0_i_s_raddr_core_sct : IN STD_LOGIC;
      twiddle_rsc_0_0_i_s_din : IN STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_s_raddr
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_s_din
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  twiddle_rsc_0_0_i : work.amba_comps.ccs_axi4_slave_mem
    GENERIC MAP(
      rscid => 0,
      depth => 64,
      op_width => 32,
      cwidth => 32,
      addr_w => 6,
      nopreload => 0,
      rst_ph => 0,
      ADDR_WIDTH => 12,
      DATA_WIDTH => 32,
      ID_WIDTH => 1,
      USER_WIDTH => 1,
      REGION_MAP_SIZE => 1,
      wBASE_ADDRESS => 0,
      rBASE_ADDRESS => 0
      )
    PORT MAP(
      ACLK => clk,
      ARESETn => '1',
      AWID => twiddle_rsc_0_0_i_AWID,
      AWADDR => twiddle_rsc_0_0_i_AWADDR,
      AWLEN => twiddle_rsc_0_0_i_AWLEN,
      AWSIZE => twiddle_rsc_0_0_i_AWSIZE,
      AWBURST => twiddle_rsc_0_0_i_AWBURST,
      AWLOCK => twiddle_rsc_0_0_AWLOCK,
      AWCACHE => twiddle_rsc_0_0_i_AWCACHE,
      AWPROT => twiddle_rsc_0_0_i_AWPROT,
      AWQOS => twiddle_rsc_0_0_i_AWQOS,
      AWREGION => twiddle_rsc_0_0_i_AWREGION,
      AWUSER => twiddle_rsc_0_0_i_AWUSER,
      AWVALID => twiddle_rsc_0_0_AWVALID,
      AWREADY => twiddle_rsc_0_0_AWREADY,
      WDATA => twiddle_rsc_0_0_i_WDATA,
      WSTRB => twiddle_rsc_0_0_i_WSTRB,
      WLAST => twiddle_rsc_0_0_WLAST,
      WUSER => twiddle_rsc_0_0_i_WUSER,
      WVALID => twiddle_rsc_0_0_WVALID,
      WREADY => twiddle_rsc_0_0_WREADY,
      BID => twiddle_rsc_0_0_i_BID,
      BRESP => twiddle_rsc_0_0_i_BRESP,
      BUSER => twiddle_rsc_0_0_i_BUSER,
      BVALID => twiddle_rsc_0_0_BVALID,
      BREADY => twiddle_rsc_0_0_BREADY,
      ARID => twiddle_rsc_0_0_i_ARID,
      ARADDR => twiddle_rsc_0_0_i_ARADDR,
      ARLEN => twiddle_rsc_0_0_i_ARLEN,
      ARSIZE => twiddle_rsc_0_0_i_ARSIZE,
      ARBURST => twiddle_rsc_0_0_i_ARBURST,
      ARLOCK => twiddle_rsc_0_0_ARLOCK,
      ARCACHE => twiddle_rsc_0_0_i_ARCACHE,
      ARPROT => twiddle_rsc_0_0_i_ARPROT,
      ARQOS => twiddle_rsc_0_0_i_ARQOS,
      ARREGION => twiddle_rsc_0_0_i_ARREGION,
      ARUSER => twiddle_rsc_0_0_i_ARUSER,
      ARVALID => twiddle_rsc_0_0_ARVALID,
      ARREADY => twiddle_rsc_0_0_ARREADY,
      RID => twiddle_rsc_0_0_i_RID,
      RDATA => twiddle_rsc_0_0_i_RDATA,
      RRESP => twiddle_rsc_0_0_i_RRESP,
      RLAST => twiddle_rsc_0_0_RLAST,
      RUSER => twiddle_rsc_0_0_i_RUSER,
      RVALID => twiddle_rsc_0_0_RVALID,
      RREADY => twiddle_rsc_0_0_RREADY,
      s_re => twiddle_rsc_0_0_i_s_re_core_sct,
      s_we => '0',
      s_raddr => twiddle_rsc_0_0_i_s_raddr_1,
      s_waddr => twiddle_rsc_0_0_i_s_waddr,
      s_din => twiddle_rsc_0_0_i_s_din_1,
      s_dout => twiddle_rsc_0_0_i_s_dout,
      s_rrdy => twiddle_rsc_0_0_i_s_rrdy,
      s_wrdy => twiddle_rsc_0_0_i_s_wrdy,
      is_idle => twiddle_rsc_0_0_is_idle,
      tr_write_done => twiddle_rsc_0_0_tr_write_done,
      s_tdone => twiddle_rsc_0_0_s_tdone
    );
  twiddle_rsc_0_0_i_AWID(0) <= twiddle_rsc_0_0_AWID;
  twiddle_rsc_0_0_i_AWADDR <= twiddle_rsc_0_0_AWADDR;
  twiddle_rsc_0_0_i_AWLEN <= twiddle_rsc_0_0_AWLEN;
  twiddle_rsc_0_0_i_AWSIZE <= twiddle_rsc_0_0_AWSIZE;
  twiddle_rsc_0_0_i_AWBURST <= twiddle_rsc_0_0_AWBURST;
  twiddle_rsc_0_0_i_AWCACHE <= twiddle_rsc_0_0_AWCACHE;
  twiddle_rsc_0_0_i_AWPROT <= twiddle_rsc_0_0_AWPROT;
  twiddle_rsc_0_0_i_AWQOS <= twiddle_rsc_0_0_AWQOS;
  twiddle_rsc_0_0_i_AWREGION <= twiddle_rsc_0_0_AWREGION;
  twiddle_rsc_0_0_i_AWUSER(0) <= twiddle_rsc_0_0_AWUSER;
  twiddle_rsc_0_0_i_WDATA <= twiddle_rsc_0_0_WDATA;
  twiddle_rsc_0_0_i_WSTRB <= twiddle_rsc_0_0_WSTRB;
  twiddle_rsc_0_0_i_WUSER(0) <= twiddle_rsc_0_0_WUSER;
  twiddle_rsc_0_0_BID <= twiddle_rsc_0_0_i_BID(0);
  twiddle_rsc_0_0_BRESP <= twiddle_rsc_0_0_i_BRESP;
  twiddle_rsc_0_0_BUSER <= twiddle_rsc_0_0_i_BUSER(0);
  twiddle_rsc_0_0_i_ARID(0) <= twiddle_rsc_0_0_ARID;
  twiddle_rsc_0_0_i_ARADDR <= twiddle_rsc_0_0_ARADDR;
  twiddle_rsc_0_0_i_ARLEN <= twiddle_rsc_0_0_ARLEN;
  twiddle_rsc_0_0_i_ARSIZE <= twiddle_rsc_0_0_ARSIZE;
  twiddle_rsc_0_0_i_ARBURST <= twiddle_rsc_0_0_ARBURST;
  twiddle_rsc_0_0_i_ARCACHE <= twiddle_rsc_0_0_ARCACHE;
  twiddle_rsc_0_0_i_ARPROT <= twiddle_rsc_0_0_ARPROT;
  twiddle_rsc_0_0_i_ARQOS <= twiddle_rsc_0_0_ARQOS;
  twiddle_rsc_0_0_i_ARREGION <= twiddle_rsc_0_0_ARREGION;
  twiddle_rsc_0_0_i_ARUSER(0) <= twiddle_rsc_0_0_ARUSER;
  twiddle_rsc_0_0_RID <= twiddle_rsc_0_0_i_RID(0);
  twiddle_rsc_0_0_RDATA <= twiddle_rsc_0_0_i_RDATA;
  twiddle_rsc_0_0_RRESP <= twiddle_rsc_0_0_i_RRESP;
  twiddle_rsc_0_0_RUSER <= twiddle_rsc_0_0_i_RUSER(0);
  twiddle_rsc_0_0_i_s_raddr_1 <= twiddle_rsc_0_0_i_s_raddr;
  twiddle_rsc_0_0_i_s_waddr <= STD_LOGIC_VECTOR'( "000000");
  twiddle_rsc_0_0_i_s_din <= twiddle_rsc_0_0_i_s_din_1;
  twiddle_rsc_0_0_i_s_dout <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");

  peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_ctrl_inst : peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      twiddle_rsc_0_0_i_oswt => twiddle_rsc_0_0_i_oswt,
      twiddle_rsc_0_0_i_biwt => twiddle_rsc_0_0_i_biwt,
      twiddle_rsc_0_0_i_bdwt => twiddle_rsc_0_0_i_bdwt,
      twiddle_rsc_0_0_i_bcwt => twiddle_rsc_0_0_i_bcwt,
      twiddle_rsc_0_0_i_s_re_core_sct => twiddle_rsc_0_0_i_s_re_core_sct,
      twiddle_rsc_0_0_i_s_rrdy => twiddle_rsc_0_0_i_s_rrdy
    );
  peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp_inst : peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_0_i_oswt => twiddle_rsc_0_0_i_oswt,
      twiddle_rsc_0_0_i_wen_comp => twiddle_rsc_0_0_i_wen_comp,
      twiddle_rsc_0_0_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_s_raddr_core,
      twiddle_rsc_0_0_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_s_din_mxwt,
      twiddle_rsc_0_0_i_biwt => twiddle_rsc_0_0_i_biwt,
      twiddle_rsc_0_0_i_bdwt => twiddle_rsc_0_0_i_bdwt,
      twiddle_rsc_0_0_i_bcwt => twiddle_rsc_0_0_i_bcwt,
      twiddle_rsc_0_0_i_s_raddr => peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_s_raddr,
      twiddle_rsc_0_0_i_s_raddr_core_sct => twiddle_rsc_0_0_i_s_re_core_sct,
      twiddle_rsc_0_0_i_s_din => peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_s_din
    );
  peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_s_raddr_core
      <= '0' & (twiddle_rsc_0_0_i_s_raddr_core(4 DOWNTO 0));
  twiddle_rsc_0_0_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_s_din_mxwt;
  twiddle_rsc_0_0_i_s_raddr <= peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_s_raddr;
  peaseNTT_core_twiddle_rsc_0_0_i_twiddle_rsc_0_0_wait_dp_inst_twiddle_rsc_0_0_i_s_din
      <= twiddle_rsc_0_0_i_s_din;

END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_31_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_31_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_31_i_oswt : IN STD_LOGIC;
    xt_rsc_1_31_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_31_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_31_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_31_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_31_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_31_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_31_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_31_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_31_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_31_i_oswt : IN STD_LOGIC;
      xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_31_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_31_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_31_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_31_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_31_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_31_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_31_i_biwt : IN STD_LOGIC;
      xt_rsc_1_31_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_dp_inst_xt_rsc_1_31_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_dp_inst_xt_rsc_1_31_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_31_i_oswt => xt_rsc_1_31_i_oswt,
      xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_31_i_biwt => xt_rsc_1_31_i_biwt,
      xt_rsc_1_31_i_bdwt => xt_rsc_1_31_i_bdwt,
      xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_31_i_wea_d_core_sct_pff => xt_rsc_1_31_i_wea_d_core_sct_iff,
      xt_rsc_1_31_i_wea_d_core_psct_pff => xt_rsc_1_31_i_wea_d_core_psct_pff,
      xt_rsc_1_31_i_oswt_pff => xt_rsc_1_31_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_dp_inst : peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_31_i_qa_d => peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_dp_inst_xt_rsc_1_31_i_qa_d,
      xt_rsc_1_31_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_dp_inst_xt_rsc_1_31_i_qa_d_mxwt,
      xt_rsc_1_31_i_biwt => xt_rsc_1_31_i_biwt,
      xt_rsc_1_31_i_bdwt => xt_rsc_1_31_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_dp_inst_xt_rsc_1_31_i_qa_d <= xt_rsc_1_31_i_qa_d;
  xt_rsc_1_31_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_31_i_1_xt_rsc_1_31_wait_dp_inst_xt_rsc_1_31_i_qa_d_mxwt;

  xt_rsc_1_31_i_wea_d_pff <= xt_rsc_1_31_i_wea_d_core_sct_iff;
  xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_30_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_30_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_30_i_oswt : IN STD_LOGIC;
    xt_rsc_1_30_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_30_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_30_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_30_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_30_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_30_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_30_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_30_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_30_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_30_i_oswt : IN STD_LOGIC;
      xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_30_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_30_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_30_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_30_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_30_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_30_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_30_i_biwt : IN STD_LOGIC;
      xt_rsc_1_30_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_dp_inst_xt_rsc_1_30_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_dp_inst_xt_rsc_1_30_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_30_i_oswt => xt_rsc_1_30_i_oswt,
      xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_30_i_biwt => xt_rsc_1_30_i_biwt,
      xt_rsc_1_30_i_bdwt => xt_rsc_1_30_i_bdwt,
      xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_30_i_wea_d_core_sct_pff => xt_rsc_1_30_i_wea_d_core_sct_iff,
      xt_rsc_1_30_i_wea_d_core_psct_pff => xt_rsc_1_30_i_wea_d_core_psct_pff,
      xt_rsc_1_30_i_oswt_pff => xt_rsc_1_30_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_dp_inst : peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_30_i_qa_d => peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_dp_inst_xt_rsc_1_30_i_qa_d,
      xt_rsc_1_30_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_dp_inst_xt_rsc_1_30_i_qa_d_mxwt,
      xt_rsc_1_30_i_biwt => xt_rsc_1_30_i_biwt,
      xt_rsc_1_30_i_bdwt => xt_rsc_1_30_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_dp_inst_xt_rsc_1_30_i_qa_d <= xt_rsc_1_30_i_qa_d;
  xt_rsc_1_30_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_30_i_1_xt_rsc_1_30_wait_dp_inst_xt_rsc_1_30_i_qa_d_mxwt;

  xt_rsc_1_30_i_wea_d_pff <= xt_rsc_1_30_i_wea_d_core_sct_iff;
  xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_29_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_29_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_29_i_oswt : IN STD_LOGIC;
    xt_rsc_1_29_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_29_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_29_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_29_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_29_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_29_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_29_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_29_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_29_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_29_i_oswt : IN STD_LOGIC;
      xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_29_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_29_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_29_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_29_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_29_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_29_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_29_i_biwt : IN STD_LOGIC;
      xt_rsc_1_29_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_dp_inst_xt_rsc_1_29_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_dp_inst_xt_rsc_1_29_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_29_i_oswt => xt_rsc_1_29_i_oswt,
      xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_29_i_biwt => xt_rsc_1_29_i_biwt,
      xt_rsc_1_29_i_bdwt => xt_rsc_1_29_i_bdwt,
      xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_29_i_wea_d_core_sct_pff => xt_rsc_1_29_i_wea_d_core_sct_iff,
      xt_rsc_1_29_i_wea_d_core_psct_pff => xt_rsc_1_29_i_wea_d_core_psct_pff,
      xt_rsc_1_29_i_oswt_pff => xt_rsc_1_29_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_dp_inst : peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_29_i_qa_d => peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_dp_inst_xt_rsc_1_29_i_qa_d,
      xt_rsc_1_29_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_dp_inst_xt_rsc_1_29_i_qa_d_mxwt,
      xt_rsc_1_29_i_biwt => xt_rsc_1_29_i_biwt,
      xt_rsc_1_29_i_bdwt => xt_rsc_1_29_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_dp_inst_xt_rsc_1_29_i_qa_d <= xt_rsc_1_29_i_qa_d;
  xt_rsc_1_29_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_29_i_1_xt_rsc_1_29_wait_dp_inst_xt_rsc_1_29_i_qa_d_mxwt;

  xt_rsc_1_29_i_wea_d_pff <= xt_rsc_1_29_i_wea_d_core_sct_iff;
  xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_28_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_28_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_28_i_oswt : IN STD_LOGIC;
    xt_rsc_1_28_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_28_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_28_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_28_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_28_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_28_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_28_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_28_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_28_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_28_i_oswt : IN STD_LOGIC;
      xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_28_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_28_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_28_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_28_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_28_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_28_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_28_i_biwt : IN STD_LOGIC;
      xt_rsc_1_28_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_dp_inst_xt_rsc_1_28_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_dp_inst_xt_rsc_1_28_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_28_i_oswt => xt_rsc_1_28_i_oswt,
      xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_28_i_biwt => xt_rsc_1_28_i_biwt,
      xt_rsc_1_28_i_bdwt => xt_rsc_1_28_i_bdwt,
      xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_28_i_wea_d_core_sct_pff => xt_rsc_1_28_i_wea_d_core_sct_iff,
      xt_rsc_1_28_i_wea_d_core_psct_pff => xt_rsc_1_28_i_wea_d_core_psct_pff,
      xt_rsc_1_28_i_oswt_pff => xt_rsc_1_28_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_dp_inst : peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_28_i_qa_d => peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_dp_inst_xt_rsc_1_28_i_qa_d,
      xt_rsc_1_28_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_dp_inst_xt_rsc_1_28_i_qa_d_mxwt,
      xt_rsc_1_28_i_biwt => xt_rsc_1_28_i_biwt,
      xt_rsc_1_28_i_bdwt => xt_rsc_1_28_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_dp_inst_xt_rsc_1_28_i_qa_d <= xt_rsc_1_28_i_qa_d;
  xt_rsc_1_28_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_28_i_1_xt_rsc_1_28_wait_dp_inst_xt_rsc_1_28_i_qa_d_mxwt;

  xt_rsc_1_28_i_wea_d_pff <= xt_rsc_1_28_i_wea_d_core_sct_iff;
  xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_27_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_27_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_27_i_oswt : IN STD_LOGIC;
    xt_rsc_1_27_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_27_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_27_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_27_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_27_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_27_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_27_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_27_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_27_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_27_i_oswt : IN STD_LOGIC;
      xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_27_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_27_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_27_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_27_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_27_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_27_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_27_i_biwt : IN STD_LOGIC;
      xt_rsc_1_27_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_dp_inst_xt_rsc_1_27_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_dp_inst_xt_rsc_1_27_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_27_i_oswt => xt_rsc_1_27_i_oswt,
      xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_27_i_biwt => xt_rsc_1_27_i_biwt,
      xt_rsc_1_27_i_bdwt => xt_rsc_1_27_i_bdwt,
      xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_27_i_wea_d_core_sct_pff => xt_rsc_1_27_i_wea_d_core_sct_iff,
      xt_rsc_1_27_i_wea_d_core_psct_pff => xt_rsc_1_27_i_wea_d_core_psct_pff,
      xt_rsc_1_27_i_oswt_pff => xt_rsc_1_27_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_dp_inst : peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_27_i_qa_d => peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_dp_inst_xt_rsc_1_27_i_qa_d,
      xt_rsc_1_27_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_dp_inst_xt_rsc_1_27_i_qa_d_mxwt,
      xt_rsc_1_27_i_biwt => xt_rsc_1_27_i_biwt,
      xt_rsc_1_27_i_bdwt => xt_rsc_1_27_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_dp_inst_xt_rsc_1_27_i_qa_d <= xt_rsc_1_27_i_qa_d;
  xt_rsc_1_27_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_27_i_1_xt_rsc_1_27_wait_dp_inst_xt_rsc_1_27_i_qa_d_mxwt;

  xt_rsc_1_27_i_wea_d_pff <= xt_rsc_1_27_i_wea_d_core_sct_iff;
  xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_26_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_26_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_26_i_oswt : IN STD_LOGIC;
    xt_rsc_1_26_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_26_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_26_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_26_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_26_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_26_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_26_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_26_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_26_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_26_i_oswt : IN STD_LOGIC;
      xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_26_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_26_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_26_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_26_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_26_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_26_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_26_i_biwt : IN STD_LOGIC;
      xt_rsc_1_26_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_dp_inst_xt_rsc_1_26_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_dp_inst_xt_rsc_1_26_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_26_i_oswt => xt_rsc_1_26_i_oswt,
      xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_26_i_biwt => xt_rsc_1_26_i_biwt,
      xt_rsc_1_26_i_bdwt => xt_rsc_1_26_i_bdwt,
      xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_26_i_wea_d_core_sct_pff => xt_rsc_1_26_i_wea_d_core_sct_iff,
      xt_rsc_1_26_i_wea_d_core_psct_pff => xt_rsc_1_26_i_wea_d_core_psct_pff,
      xt_rsc_1_26_i_oswt_pff => xt_rsc_1_26_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_dp_inst : peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_26_i_qa_d => peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_dp_inst_xt_rsc_1_26_i_qa_d,
      xt_rsc_1_26_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_dp_inst_xt_rsc_1_26_i_qa_d_mxwt,
      xt_rsc_1_26_i_biwt => xt_rsc_1_26_i_biwt,
      xt_rsc_1_26_i_bdwt => xt_rsc_1_26_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_dp_inst_xt_rsc_1_26_i_qa_d <= xt_rsc_1_26_i_qa_d;
  xt_rsc_1_26_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_26_i_1_xt_rsc_1_26_wait_dp_inst_xt_rsc_1_26_i_qa_d_mxwt;

  xt_rsc_1_26_i_wea_d_pff <= xt_rsc_1_26_i_wea_d_core_sct_iff;
  xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_25_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_25_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_25_i_oswt : IN STD_LOGIC;
    xt_rsc_1_25_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_25_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_25_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_25_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_25_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_25_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_25_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_25_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_25_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_25_i_oswt : IN STD_LOGIC;
      xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_25_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_25_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_25_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_25_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_25_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_25_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_25_i_biwt : IN STD_LOGIC;
      xt_rsc_1_25_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_dp_inst_xt_rsc_1_25_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_dp_inst_xt_rsc_1_25_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_25_i_oswt => xt_rsc_1_25_i_oswt,
      xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_25_i_biwt => xt_rsc_1_25_i_biwt,
      xt_rsc_1_25_i_bdwt => xt_rsc_1_25_i_bdwt,
      xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_25_i_wea_d_core_sct_pff => xt_rsc_1_25_i_wea_d_core_sct_iff,
      xt_rsc_1_25_i_wea_d_core_psct_pff => xt_rsc_1_25_i_wea_d_core_psct_pff,
      xt_rsc_1_25_i_oswt_pff => xt_rsc_1_25_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_dp_inst : peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_25_i_qa_d => peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_dp_inst_xt_rsc_1_25_i_qa_d,
      xt_rsc_1_25_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_dp_inst_xt_rsc_1_25_i_qa_d_mxwt,
      xt_rsc_1_25_i_biwt => xt_rsc_1_25_i_biwt,
      xt_rsc_1_25_i_bdwt => xt_rsc_1_25_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_dp_inst_xt_rsc_1_25_i_qa_d <= xt_rsc_1_25_i_qa_d;
  xt_rsc_1_25_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_25_i_1_xt_rsc_1_25_wait_dp_inst_xt_rsc_1_25_i_qa_d_mxwt;

  xt_rsc_1_25_i_wea_d_pff <= xt_rsc_1_25_i_wea_d_core_sct_iff;
  xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_24_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_24_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_24_i_oswt : IN STD_LOGIC;
    xt_rsc_1_24_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_24_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_24_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_24_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_24_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_24_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_24_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_24_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_24_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_24_i_oswt : IN STD_LOGIC;
      xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_24_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_24_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_24_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_24_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_24_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_24_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_24_i_biwt : IN STD_LOGIC;
      xt_rsc_1_24_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_dp_inst_xt_rsc_1_24_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_dp_inst_xt_rsc_1_24_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_24_i_oswt => xt_rsc_1_24_i_oswt,
      xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_24_i_biwt => xt_rsc_1_24_i_biwt,
      xt_rsc_1_24_i_bdwt => xt_rsc_1_24_i_bdwt,
      xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_24_i_wea_d_core_sct_pff => xt_rsc_1_24_i_wea_d_core_sct_iff,
      xt_rsc_1_24_i_wea_d_core_psct_pff => xt_rsc_1_24_i_wea_d_core_psct_pff,
      xt_rsc_1_24_i_oswt_pff => xt_rsc_1_24_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_dp_inst : peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_24_i_qa_d => peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_dp_inst_xt_rsc_1_24_i_qa_d,
      xt_rsc_1_24_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_dp_inst_xt_rsc_1_24_i_qa_d_mxwt,
      xt_rsc_1_24_i_biwt => xt_rsc_1_24_i_biwt,
      xt_rsc_1_24_i_bdwt => xt_rsc_1_24_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_dp_inst_xt_rsc_1_24_i_qa_d <= xt_rsc_1_24_i_qa_d;
  xt_rsc_1_24_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_24_i_1_xt_rsc_1_24_wait_dp_inst_xt_rsc_1_24_i_qa_d_mxwt;

  xt_rsc_1_24_i_wea_d_pff <= xt_rsc_1_24_i_wea_d_core_sct_iff;
  xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_23_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_23_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_23_i_oswt : IN STD_LOGIC;
    xt_rsc_1_23_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_23_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_23_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_23_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_23_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_23_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_23_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_23_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_23_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_23_i_oswt : IN STD_LOGIC;
      xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_23_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_23_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_23_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_23_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_23_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_23_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_23_i_biwt : IN STD_LOGIC;
      xt_rsc_1_23_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_dp_inst_xt_rsc_1_23_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_dp_inst_xt_rsc_1_23_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_23_i_oswt => xt_rsc_1_23_i_oswt,
      xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_23_i_biwt => xt_rsc_1_23_i_biwt,
      xt_rsc_1_23_i_bdwt => xt_rsc_1_23_i_bdwt,
      xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_23_i_wea_d_core_sct_pff => xt_rsc_1_23_i_wea_d_core_sct_iff,
      xt_rsc_1_23_i_wea_d_core_psct_pff => xt_rsc_1_23_i_wea_d_core_psct_pff,
      xt_rsc_1_23_i_oswt_pff => xt_rsc_1_23_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_dp_inst : peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_23_i_qa_d => peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_dp_inst_xt_rsc_1_23_i_qa_d,
      xt_rsc_1_23_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_dp_inst_xt_rsc_1_23_i_qa_d_mxwt,
      xt_rsc_1_23_i_biwt => xt_rsc_1_23_i_biwt,
      xt_rsc_1_23_i_bdwt => xt_rsc_1_23_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_dp_inst_xt_rsc_1_23_i_qa_d <= xt_rsc_1_23_i_qa_d;
  xt_rsc_1_23_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_23_i_1_xt_rsc_1_23_wait_dp_inst_xt_rsc_1_23_i_qa_d_mxwt;

  xt_rsc_1_23_i_wea_d_pff <= xt_rsc_1_23_i_wea_d_core_sct_iff;
  xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_22_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_22_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_22_i_oswt : IN STD_LOGIC;
    xt_rsc_1_22_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_22_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_22_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_22_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_22_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_22_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_22_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_22_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_22_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_22_i_oswt : IN STD_LOGIC;
      xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_22_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_22_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_22_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_22_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_22_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_22_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_22_i_biwt : IN STD_LOGIC;
      xt_rsc_1_22_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_dp_inst_xt_rsc_1_22_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_dp_inst_xt_rsc_1_22_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_22_i_oswt => xt_rsc_1_22_i_oswt,
      xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_22_i_biwt => xt_rsc_1_22_i_biwt,
      xt_rsc_1_22_i_bdwt => xt_rsc_1_22_i_bdwt,
      xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_22_i_wea_d_core_sct_pff => xt_rsc_1_22_i_wea_d_core_sct_iff,
      xt_rsc_1_22_i_wea_d_core_psct_pff => xt_rsc_1_22_i_wea_d_core_psct_pff,
      xt_rsc_1_22_i_oswt_pff => xt_rsc_1_22_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_dp_inst : peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_22_i_qa_d => peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_dp_inst_xt_rsc_1_22_i_qa_d,
      xt_rsc_1_22_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_dp_inst_xt_rsc_1_22_i_qa_d_mxwt,
      xt_rsc_1_22_i_biwt => xt_rsc_1_22_i_biwt,
      xt_rsc_1_22_i_bdwt => xt_rsc_1_22_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_dp_inst_xt_rsc_1_22_i_qa_d <= xt_rsc_1_22_i_qa_d;
  xt_rsc_1_22_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_22_i_1_xt_rsc_1_22_wait_dp_inst_xt_rsc_1_22_i_qa_d_mxwt;

  xt_rsc_1_22_i_wea_d_pff <= xt_rsc_1_22_i_wea_d_core_sct_iff;
  xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_21_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_21_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_21_i_oswt : IN STD_LOGIC;
    xt_rsc_1_21_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_21_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_21_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_21_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_21_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_21_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_21_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_21_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_21_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_21_i_oswt : IN STD_LOGIC;
      xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_21_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_21_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_21_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_21_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_21_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_21_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_21_i_biwt : IN STD_LOGIC;
      xt_rsc_1_21_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_dp_inst_xt_rsc_1_21_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_dp_inst_xt_rsc_1_21_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_21_i_oswt => xt_rsc_1_21_i_oswt,
      xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_21_i_biwt => xt_rsc_1_21_i_biwt,
      xt_rsc_1_21_i_bdwt => xt_rsc_1_21_i_bdwt,
      xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_21_i_wea_d_core_sct_pff => xt_rsc_1_21_i_wea_d_core_sct_iff,
      xt_rsc_1_21_i_wea_d_core_psct_pff => xt_rsc_1_21_i_wea_d_core_psct_pff,
      xt_rsc_1_21_i_oswt_pff => xt_rsc_1_21_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_dp_inst : peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_21_i_qa_d => peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_dp_inst_xt_rsc_1_21_i_qa_d,
      xt_rsc_1_21_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_dp_inst_xt_rsc_1_21_i_qa_d_mxwt,
      xt_rsc_1_21_i_biwt => xt_rsc_1_21_i_biwt,
      xt_rsc_1_21_i_bdwt => xt_rsc_1_21_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_dp_inst_xt_rsc_1_21_i_qa_d <= xt_rsc_1_21_i_qa_d;
  xt_rsc_1_21_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_21_i_1_xt_rsc_1_21_wait_dp_inst_xt_rsc_1_21_i_qa_d_mxwt;

  xt_rsc_1_21_i_wea_d_pff <= xt_rsc_1_21_i_wea_d_core_sct_iff;
  xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_20_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_20_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_20_i_oswt : IN STD_LOGIC;
    xt_rsc_1_20_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_20_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_20_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_20_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_20_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_20_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_20_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_20_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_20_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_20_i_oswt : IN STD_LOGIC;
      xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_20_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_20_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_20_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_20_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_20_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_20_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_20_i_biwt : IN STD_LOGIC;
      xt_rsc_1_20_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_dp_inst_xt_rsc_1_20_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_dp_inst_xt_rsc_1_20_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_20_i_oswt => xt_rsc_1_20_i_oswt,
      xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_20_i_biwt => xt_rsc_1_20_i_biwt,
      xt_rsc_1_20_i_bdwt => xt_rsc_1_20_i_bdwt,
      xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_20_i_wea_d_core_sct_pff => xt_rsc_1_20_i_wea_d_core_sct_iff,
      xt_rsc_1_20_i_wea_d_core_psct_pff => xt_rsc_1_20_i_wea_d_core_psct_pff,
      xt_rsc_1_20_i_oswt_pff => xt_rsc_1_20_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_dp_inst : peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_20_i_qa_d => peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_dp_inst_xt_rsc_1_20_i_qa_d,
      xt_rsc_1_20_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_dp_inst_xt_rsc_1_20_i_qa_d_mxwt,
      xt_rsc_1_20_i_biwt => xt_rsc_1_20_i_biwt,
      xt_rsc_1_20_i_bdwt => xt_rsc_1_20_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_dp_inst_xt_rsc_1_20_i_qa_d <= xt_rsc_1_20_i_qa_d;
  xt_rsc_1_20_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_20_i_1_xt_rsc_1_20_wait_dp_inst_xt_rsc_1_20_i_qa_d_mxwt;

  xt_rsc_1_20_i_wea_d_pff <= xt_rsc_1_20_i_wea_d_core_sct_iff;
  xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_19_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_19_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_19_i_oswt : IN STD_LOGIC;
    xt_rsc_1_19_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_19_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_19_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_19_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_19_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_19_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_19_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_19_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_19_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_19_i_oswt : IN STD_LOGIC;
      xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_19_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_19_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_19_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_19_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_19_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_19_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_19_i_biwt : IN STD_LOGIC;
      xt_rsc_1_19_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_dp_inst_xt_rsc_1_19_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_dp_inst_xt_rsc_1_19_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_19_i_oswt => xt_rsc_1_19_i_oswt,
      xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_19_i_biwt => xt_rsc_1_19_i_biwt,
      xt_rsc_1_19_i_bdwt => xt_rsc_1_19_i_bdwt,
      xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_19_i_wea_d_core_sct_pff => xt_rsc_1_19_i_wea_d_core_sct_iff,
      xt_rsc_1_19_i_wea_d_core_psct_pff => xt_rsc_1_19_i_wea_d_core_psct_pff,
      xt_rsc_1_19_i_oswt_pff => xt_rsc_1_19_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_dp_inst : peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_19_i_qa_d => peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_dp_inst_xt_rsc_1_19_i_qa_d,
      xt_rsc_1_19_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_dp_inst_xt_rsc_1_19_i_qa_d_mxwt,
      xt_rsc_1_19_i_biwt => xt_rsc_1_19_i_biwt,
      xt_rsc_1_19_i_bdwt => xt_rsc_1_19_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_dp_inst_xt_rsc_1_19_i_qa_d <= xt_rsc_1_19_i_qa_d;
  xt_rsc_1_19_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_19_i_1_xt_rsc_1_19_wait_dp_inst_xt_rsc_1_19_i_qa_d_mxwt;

  xt_rsc_1_19_i_wea_d_pff <= xt_rsc_1_19_i_wea_d_core_sct_iff;
  xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_18_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_18_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_18_i_oswt : IN STD_LOGIC;
    xt_rsc_1_18_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_18_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_18_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_18_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_18_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_18_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_18_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_18_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_18_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_18_i_oswt : IN STD_LOGIC;
      xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_18_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_18_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_18_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_18_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_18_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_18_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_18_i_biwt : IN STD_LOGIC;
      xt_rsc_1_18_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_dp_inst_xt_rsc_1_18_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_dp_inst_xt_rsc_1_18_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_18_i_oswt => xt_rsc_1_18_i_oswt,
      xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_18_i_biwt => xt_rsc_1_18_i_biwt,
      xt_rsc_1_18_i_bdwt => xt_rsc_1_18_i_bdwt,
      xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_18_i_wea_d_core_sct_pff => xt_rsc_1_18_i_wea_d_core_sct_iff,
      xt_rsc_1_18_i_wea_d_core_psct_pff => xt_rsc_1_18_i_wea_d_core_psct_pff,
      xt_rsc_1_18_i_oswt_pff => xt_rsc_1_18_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_dp_inst : peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_18_i_qa_d => peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_dp_inst_xt_rsc_1_18_i_qa_d,
      xt_rsc_1_18_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_dp_inst_xt_rsc_1_18_i_qa_d_mxwt,
      xt_rsc_1_18_i_biwt => xt_rsc_1_18_i_biwt,
      xt_rsc_1_18_i_bdwt => xt_rsc_1_18_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_dp_inst_xt_rsc_1_18_i_qa_d <= xt_rsc_1_18_i_qa_d;
  xt_rsc_1_18_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_18_i_1_xt_rsc_1_18_wait_dp_inst_xt_rsc_1_18_i_qa_d_mxwt;

  xt_rsc_1_18_i_wea_d_pff <= xt_rsc_1_18_i_wea_d_core_sct_iff;
  xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_17_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_17_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_17_i_oswt : IN STD_LOGIC;
    xt_rsc_1_17_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_17_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_17_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_17_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_17_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_17_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_17_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_17_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_17_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_17_i_oswt : IN STD_LOGIC;
      xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_17_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_17_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_17_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_17_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_17_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_17_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_17_i_biwt : IN STD_LOGIC;
      xt_rsc_1_17_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_dp_inst_xt_rsc_1_17_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_dp_inst_xt_rsc_1_17_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_17_i_oswt => xt_rsc_1_17_i_oswt,
      xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_17_i_biwt => xt_rsc_1_17_i_biwt,
      xt_rsc_1_17_i_bdwt => xt_rsc_1_17_i_bdwt,
      xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_17_i_wea_d_core_sct_pff => xt_rsc_1_17_i_wea_d_core_sct_iff,
      xt_rsc_1_17_i_wea_d_core_psct_pff => xt_rsc_1_17_i_wea_d_core_psct_pff,
      xt_rsc_1_17_i_oswt_pff => xt_rsc_1_17_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_dp_inst : peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_17_i_qa_d => peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_dp_inst_xt_rsc_1_17_i_qa_d,
      xt_rsc_1_17_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_dp_inst_xt_rsc_1_17_i_qa_d_mxwt,
      xt_rsc_1_17_i_biwt => xt_rsc_1_17_i_biwt,
      xt_rsc_1_17_i_bdwt => xt_rsc_1_17_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_dp_inst_xt_rsc_1_17_i_qa_d <= xt_rsc_1_17_i_qa_d;
  xt_rsc_1_17_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_17_i_1_xt_rsc_1_17_wait_dp_inst_xt_rsc_1_17_i_qa_d_mxwt;

  xt_rsc_1_17_i_wea_d_pff <= xt_rsc_1_17_i_wea_d_core_sct_iff;
  xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_16_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_16_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_16_i_oswt : IN STD_LOGIC;
    xt_rsc_1_16_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_16_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_16_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_16_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_16_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_16_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_16_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_16_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_16_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_16_i_oswt : IN STD_LOGIC;
      xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_16_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_16_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_16_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_16_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_16_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_16_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_16_i_biwt : IN STD_LOGIC;
      xt_rsc_1_16_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_dp_inst_xt_rsc_1_16_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_dp_inst_xt_rsc_1_16_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_16_i_oswt => xt_rsc_1_16_i_oswt,
      xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_16_i_biwt => xt_rsc_1_16_i_biwt,
      xt_rsc_1_16_i_bdwt => xt_rsc_1_16_i_bdwt,
      xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_16_i_wea_d_core_sct_pff => xt_rsc_1_16_i_wea_d_core_sct_iff,
      xt_rsc_1_16_i_wea_d_core_psct_pff => xt_rsc_1_16_i_wea_d_core_psct_pff,
      xt_rsc_1_16_i_oswt_pff => xt_rsc_1_16_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_dp_inst : peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_16_i_qa_d => peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_dp_inst_xt_rsc_1_16_i_qa_d,
      xt_rsc_1_16_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_dp_inst_xt_rsc_1_16_i_qa_d_mxwt,
      xt_rsc_1_16_i_biwt => xt_rsc_1_16_i_biwt,
      xt_rsc_1_16_i_bdwt => xt_rsc_1_16_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_dp_inst_xt_rsc_1_16_i_qa_d <= xt_rsc_1_16_i_qa_d;
  xt_rsc_1_16_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_16_i_1_xt_rsc_1_16_wait_dp_inst_xt_rsc_1_16_i_qa_d_mxwt;

  xt_rsc_1_16_i_wea_d_pff <= xt_rsc_1_16_i_wea_d_core_sct_iff;
  xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_15_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_15_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_15_i_oswt : IN STD_LOGIC;
    xt_rsc_1_15_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_15_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_15_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_15_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_15_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_15_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_15_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_15_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_15_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_15_i_oswt : IN STD_LOGIC;
      xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_15_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_15_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_15_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_15_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_15_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_15_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_15_i_biwt : IN STD_LOGIC;
      xt_rsc_1_15_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_dp_inst_xt_rsc_1_15_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_dp_inst_xt_rsc_1_15_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_15_i_oswt => xt_rsc_1_15_i_oswt,
      xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_15_i_biwt => xt_rsc_1_15_i_biwt,
      xt_rsc_1_15_i_bdwt => xt_rsc_1_15_i_bdwt,
      xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_15_i_wea_d_core_sct_pff => xt_rsc_1_15_i_wea_d_core_sct_iff,
      xt_rsc_1_15_i_wea_d_core_psct_pff => xt_rsc_1_15_i_wea_d_core_psct_pff,
      xt_rsc_1_15_i_oswt_pff => xt_rsc_1_15_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_dp_inst : peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_15_i_qa_d => peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_dp_inst_xt_rsc_1_15_i_qa_d,
      xt_rsc_1_15_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_dp_inst_xt_rsc_1_15_i_qa_d_mxwt,
      xt_rsc_1_15_i_biwt => xt_rsc_1_15_i_biwt,
      xt_rsc_1_15_i_bdwt => xt_rsc_1_15_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_dp_inst_xt_rsc_1_15_i_qa_d <= xt_rsc_1_15_i_qa_d;
  xt_rsc_1_15_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_15_i_1_xt_rsc_1_15_wait_dp_inst_xt_rsc_1_15_i_qa_d_mxwt;

  xt_rsc_1_15_i_wea_d_pff <= xt_rsc_1_15_i_wea_d_core_sct_iff;
  xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_14_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_14_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_14_i_oswt : IN STD_LOGIC;
    xt_rsc_1_14_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_14_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_14_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_14_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_14_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_14_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_14_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_14_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_14_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_14_i_oswt : IN STD_LOGIC;
      xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_14_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_14_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_14_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_14_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_14_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_14_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_14_i_biwt : IN STD_LOGIC;
      xt_rsc_1_14_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_dp_inst_xt_rsc_1_14_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_dp_inst_xt_rsc_1_14_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_14_i_oswt => xt_rsc_1_14_i_oswt,
      xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_14_i_biwt => xt_rsc_1_14_i_biwt,
      xt_rsc_1_14_i_bdwt => xt_rsc_1_14_i_bdwt,
      xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_14_i_wea_d_core_sct_pff => xt_rsc_1_14_i_wea_d_core_sct_iff,
      xt_rsc_1_14_i_wea_d_core_psct_pff => xt_rsc_1_14_i_wea_d_core_psct_pff,
      xt_rsc_1_14_i_oswt_pff => xt_rsc_1_14_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_dp_inst : peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_14_i_qa_d => peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_dp_inst_xt_rsc_1_14_i_qa_d,
      xt_rsc_1_14_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_dp_inst_xt_rsc_1_14_i_qa_d_mxwt,
      xt_rsc_1_14_i_biwt => xt_rsc_1_14_i_biwt,
      xt_rsc_1_14_i_bdwt => xt_rsc_1_14_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_dp_inst_xt_rsc_1_14_i_qa_d <= xt_rsc_1_14_i_qa_d;
  xt_rsc_1_14_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_14_i_1_xt_rsc_1_14_wait_dp_inst_xt_rsc_1_14_i_qa_d_mxwt;

  xt_rsc_1_14_i_wea_d_pff <= xt_rsc_1_14_i_wea_d_core_sct_iff;
  xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_13_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_13_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_13_i_oswt : IN STD_LOGIC;
    xt_rsc_1_13_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_13_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_13_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_13_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_13_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_13_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_13_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_13_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_13_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_13_i_oswt : IN STD_LOGIC;
      xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_13_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_13_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_13_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_13_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_13_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_13_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_13_i_biwt : IN STD_LOGIC;
      xt_rsc_1_13_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_dp_inst_xt_rsc_1_13_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_dp_inst_xt_rsc_1_13_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_13_i_oswt => xt_rsc_1_13_i_oswt,
      xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_13_i_biwt => xt_rsc_1_13_i_biwt,
      xt_rsc_1_13_i_bdwt => xt_rsc_1_13_i_bdwt,
      xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_13_i_wea_d_core_sct_pff => xt_rsc_1_13_i_wea_d_core_sct_iff,
      xt_rsc_1_13_i_wea_d_core_psct_pff => xt_rsc_1_13_i_wea_d_core_psct_pff,
      xt_rsc_1_13_i_oswt_pff => xt_rsc_1_13_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_dp_inst : peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_13_i_qa_d => peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_dp_inst_xt_rsc_1_13_i_qa_d,
      xt_rsc_1_13_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_dp_inst_xt_rsc_1_13_i_qa_d_mxwt,
      xt_rsc_1_13_i_biwt => xt_rsc_1_13_i_biwt,
      xt_rsc_1_13_i_bdwt => xt_rsc_1_13_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_dp_inst_xt_rsc_1_13_i_qa_d <= xt_rsc_1_13_i_qa_d;
  xt_rsc_1_13_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_13_i_1_xt_rsc_1_13_wait_dp_inst_xt_rsc_1_13_i_qa_d_mxwt;

  xt_rsc_1_13_i_wea_d_pff <= xt_rsc_1_13_i_wea_d_core_sct_iff;
  xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_12_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_12_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_12_i_oswt : IN STD_LOGIC;
    xt_rsc_1_12_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_12_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_12_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_12_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_12_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_12_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_12_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_12_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_12_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_12_i_oswt : IN STD_LOGIC;
      xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_12_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_12_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_12_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_12_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_12_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_12_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_12_i_biwt : IN STD_LOGIC;
      xt_rsc_1_12_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_dp_inst_xt_rsc_1_12_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_dp_inst_xt_rsc_1_12_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_12_i_oswt => xt_rsc_1_12_i_oswt,
      xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_12_i_biwt => xt_rsc_1_12_i_biwt,
      xt_rsc_1_12_i_bdwt => xt_rsc_1_12_i_bdwt,
      xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_12_i_wea_d_core_sct_pff => xt_rsc_1_12_i_wea_d_core_sct_iff,
      xt_rsc_1_12_i_wea_d_core_psct_pff => xt_rsc_1_12_i_wea_d_core_psct_pff,
      xt_rsc_1_12_i_oswt_pff => xt_rsc_1_12_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_dp_inst : peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_12_i_qa_d => peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_dp_inst_xt_rsc_1_12_i_qa_d,
      xt_rsc_1_12_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_dp_inst_xt_rsc_1_12_i_qa_d_mxwt,
      xt_rsc_1_12_i_biwt => xt_rsc_1_12_i_biwt,
      xt_rsc_1_12_i_bdwt => xt_rsc_1_12_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_dp_inst_xt_rsc_1_12_i_qa_d <= xt_rsc_1_12_i_qa_d;
  xt_rsc_1_12_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_12_i_1_xt_rsc_1_12_wait_dp_inst_xt_rsc_1_12_i_qa_d_mxwt;

  xt_rsc_1_12_i_wea_d_pff <= xt_rsc_1_12_i_wea_d_core_sct_iff;
  xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_11_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_11_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_11_i_oswt : IN STD_LOGIC;
    xt_rsc_1_11_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_11_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_11_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_11_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_11_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_11_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_11_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_11_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_11_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_11_i_oswt : IN STD_LOGIC;
      xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_11_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_11_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_11_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_11_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_11_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_11_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_11_i_biwt : IN STD_LOGIC;
      xt_rsc_1_11_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_dp_inst_xt_rsc_1_11_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_dp_inst_xt_rsc_1_11_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_11_i_oswt => xt_rsc_1_11_i_oswt,
      xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_11_i_biwt => xt_rsc_1_11_i_biwt,
      xt_rsc_1_11_i_bdwt => xt_rsc_1_11_i_bdwt,
      xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_11_i_wea_d_core_sct_pff => xt_rsc_1_11_i_wea_d_core_sct_iff,
      xt_rsc_1_11_i_wea_d_core_psct_pff => xt_rsc_1_11_i_wea_d_core_psct_pff,
      xt_rsc_1_11_i_oswt_pff => xt_rsc_1_11_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_dp_inst : peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_11_i_qa_d => peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_dp_inst_xt_rsc_1_11_i_qa_d,
      xt_rsc_1_11_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_dp_inst_xt_rsc_1_11_i_qa_d_mxwt,
      xt_rsc_1_11_i_biwt => xt_rsc_1_11_i_biwt,
      xt_rsc_1_11_i_bdwt => xt_rsc_1_11_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_dp_inst_xt_rsc_1_11_i_qa_d <= xt_rsc_1_11_i_qa_d;
  xt_rsc_1_11_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_11_i_1_xt_rsc_1_11_wait_dp_inst_xt_rsc_1_11_i_qa_d_mxwt;

  xt_rsc_1_11_i_wea_d_pff <= xt_rsc_1_11_i_wea_d_core_sct_iff;
  xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_10_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_10_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_10_i_oswt : IN STD_LOGIC;
    xt_rsc_1_10_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_10_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_10_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_10_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_10_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_10_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_10_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_10_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_10_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_10_i_oswt : IN STD_LOGIC;
      xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_10_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_10_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_10_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_10_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_10_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_10_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_10_i_biwt : IN STD_LOGIC;
      xt_rsc_1_10_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_dp_inst_xt_rsc_1_10_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_dp_inst_xt_rsc_1_10_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_10_i_oswt => xt_rsc_1_10_i_oswt,
      xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_10_i_biwt => xt_rsc_1_10_i_biwt,
      xt_rsc_1_10_i_bdwt => xt_rsc_1_10_i_bdwt,
      xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_10_i_wea_d_core_sct_pff => xt_rsc_1_10_i_wea_d_core_sct_iff,
      xt_rsc_1_10_i_wea_d_core_psct_pff => xt_rsc_1_10_i_wea_d_core_psct_pff,
      xt_rsc_1_10_i_oswt_pff => xt_rsc_1_10_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_dp_inst : peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_10_i_qa_d => peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_dp_inst_xt_rsc_1_10_i_qa_d,
      xt_rsc_1_10_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_dp_inst_xt_rsc_1_10_i_qa_d_mxwt,
      xt_rsc_1_10_i_biwt => xt_rsc_1_10_i_biwt,
      xt_rsc_1_10_i_bdwt => xt_rsc_1_10_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_dp_inst_xt_rsc_1_10_i_qa_d <= xt_rsc_1_10_i_qa_d;
  xt_rsc_1_10_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_10_i_1_xt_rsc_1_10_wait_dp_inst_xt_rsc_1_10_i_qa_d_mxwt;

  xt_rsc_1_10_i_wea_d_pff <= xt_rsc_1_10_i_wea_d_core_sct_iff;
  xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_9_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_9_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_9_i_oswt : IN STD_LOGIC;
    xt_rsc_1_9_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_9_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_9_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_9_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_9_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_9_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_9_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_9_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_9_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_9_i_oswt : IN STD_LOGIC;
      xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_9_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_9_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_9_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_9_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_9_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_9_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_9_i_biwt : IN STD_LOGIC;
      xt_rsc_1_9_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_dp_inst_xt_rsc_1_9_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_dp_inst_xt_rsc_1_9_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_9_i_oswt => xt_rsc_1_9_i_oswt,
      xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_9_i_biwt => xt_rsc_1_9_i_biwt,
      xt_rsc_1_9_i_bdwt => xt_rsc_1_9_i_bdwt,
      xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_9_i_wea_d_core_sct_pff => xt_rsc_1_9_i_wea_d_core_sct_iff,
      xt_rsc_1_9_i_wea_d_core_psct_pff => xt_rsc_1_9_i_wea_d_core_psct_pff,
      xt_rsc_1_9_i_oswt_pff => xt_rsc_1_9_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_dp_inst : peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_9_i_qa_d => peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_dp_inst_xt_rsc_1_9_i_qa_d,
      xt_rsc_1_9_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_dp_inst_xt_rsc_1_9_i_qa_d_mxwt,
      xt_rsc_1_9_i_biwt => xt_rsc_1_9_i_biwt,
      xt_rsc_1_9_i_bdwt => xt_rsc_1_9_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_dp_inst_xt_rsc_1_9_i_qa_d <= xt_rsc_1_9_i_qa_d;
  xt_rsc_1_9_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_9_i_1_xt_rsc_1_9_wait_dp_inst_xt_rsc_1_9_i_qa_d_mxwt;

  xt_rsc_1_9_i_wea_d_pff <= xt_rsc_1_9_i_wea_d_core_sct_iff;
  xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_8_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_8_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_8_i_oswt : IN STD_LOGIC;
    xt_rsc_1_8_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_8_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_8_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_8_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_8_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_8_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_8_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_8_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_8_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_8_i_oswt : IN STD_LOGIC;
      xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_8_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_8_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_8_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_8_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_8_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_8_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_8_i_biwt : IN STD_LOGIC;
      xt_rsc_1_8_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_dp_inst_xt_rsc_1_8_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_dp_inst_xt_rsc_1_8_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_8_i_oswt => xt_rsc_1_8_i_oswt,
      xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_8_i_biwt => xt_rsc_1_8_i_biwt,
      xt_rsc_1_8_i_bdwt => xt_rsc_1_8_i_bdwt,
      xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_8_i_wea_d_core_sct_pff => xt_rsc_1_8_i_wea_d_core_sct_iff,
      xt_rsc_1_8_i_wea_d_core_psct_pff => xt_rsc_1_8_i_wea_d_core_psct_pff,
      xt_rsc_1_8_i_oswt_pff => xt_rsc_1_8_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_dp_inst : peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_8_i_qa_d => peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_dp_inst_xt_rsc_1_8_i_qa_d,
      xt_rsc_1_8_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_dp_inst_xt_rsc_1_8_i_qa_d_mxwt,
      xt_rsc_1_8_i_biwt => xt_rsc_1_8_i_biwt,
      xt_rsc_1_8_i_bdwt => xt_rsc_1_8_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_dp_inst_xt_rsc_1_8_i_qa_d <= xt_rsc_1_8_i_qa_d;
  xt_rsc_1_8_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_8_i_1_xt_rsc_1_8_wait_dp_inst_xt_rsc_1_8_i_qa_d_mxwt;

  xt_rsc_1_8_i_wea_d_pff <= xt_rsc_1_8_i_wea_d_core_sct_iff;
  xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_7_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_7_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_7_i_oswt : IN STD_LOGIC;
    xt_rsc_1_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_7_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_7_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_7_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_7_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_7_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_7_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_7_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_7_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_7_i_oswt : IN STD_LOGIC;
      xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_7_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_7_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_7_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_7_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_7_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_7_i_biwt : IN STD_LOGIC;
      xt_rsc_1_7_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_dp_inst_xt_rsc_1_7_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_dp_inst_xt_rsc_1_7_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_7_i_oswt => xt_rsc_1_7_i_oswt,
      xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_7_i_biwt => xt_rsc_1_7_i_biwt,
      xt_rsc_1_7_i_bdwt => xt_rsc_1_7_i_bdwt,
      xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_7_i_wea_d_core_sct_pff => xt_rsc_1_7_i_wea_d_core_sct_iff,
      xt_rsc_1_7_i_wea_d_core_psct_pff => xt_rsc_1_7_i_wea_d_core_psct_pff,
      xt_rsc_1_7_i_oswt_pff => xt_rsc_1_7_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_dp_inst : peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_7_i_qa_d => peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_dp_inst_xt_rsc_1_7_i_qa_d,
      xt_rsc_1_7_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_dp_inst_xt_rsc_1_7_i_qa_d_mxwt,
      xt_rsc_1_7_i_biwt => xt_rsc_1_7_i_biwt,
      xt_rsc_1_7_i_bdwt => xt_rsc_1_7_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_dp_inst_xt_rsc_1_7_i_qa_d <= xt_rsc_1_7_i_qa_d;
  xt_rsc_1_7_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_7_i_1_xt_rsc_1_7_wait_dp_inst_xt_rsc_1_7_i_qa_d_mxwt;

  xt_rsc_1_7_i_wea_d_pff <= xt_rsc_1_7_i_wea_d_core_sct_iff;
  xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_6_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_6_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_6_i_oswt : IN STD_LOGIC;
    xt_rsc_1_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_6_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_6_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_6_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_6_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_6_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_6_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_6_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_6_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_6_i_oswt : IN STD_LOGIC;
      xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_6_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_6_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_6_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_6_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_6_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_6_i_biwt : IN STD_LOGIC;
      xt_rsc_1_6_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_dp_inst_xt_rsc_1_6_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_dp_inst_xt_rsc_1_6_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_6_i_oswt => xt_rsc_1_6_i_oswt,
      xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_6_i_biwt => xt_rsc_1_6_i_biwt,
      xt_rsc_1_6_i_bdwt => xt_rsc_1_6_i_bdwt,
      xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_6_i_wea_d_core_sct_pff => xt_rsc_1_6_i_wea_d_core_sct_iff,
      xt_rsc_1_6_i_wea_d_core_psct_pff => xt_rsc_1_6_i_wea_d_core_psct_pff,
      xt_rsc_1_6_i_oswt_pff => xt_rsc_1_6_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_dp_inst : peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_6_i_qa_d => peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_dp_inst_xt_rsc_1_6_i_qa_d,
      xt_rsc_1_6_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_dp_inst_xt_rsc_1_6_i_qa_d_mxwt,
      xt_rsc_1_6_i_biwt => xt_rsc_1_6_i_biwt,
      xt_rsc_1_6_i_bdwt => xt_rsc_1_6_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_dp_inst_xt_rsc_1_6_i_qa_d <= xt_rsc_1_6_i_qa_d;
  xt_rsc_1_6_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_6_i_1_xt_rsc_1_6_wait_dp_inst_xt_rsc_1_6_i_qa_d_mxwt;

  xt_rsc_1_6_i_wea_d_pff <= xt_rsc_1_6_i_wea_d_core_sct_iff;
  xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_5_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_5_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_5_i_oswt : IN STD_LOGIC;
    xt_rsc_1_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_5_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_5_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_5_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_5_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_5_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_5_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_5_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_5_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_5_i_oswt : IN STD_LOGIC;
      xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_5_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_5_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_5_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_5_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_5_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_5_i_biwt : IN STD_LOGIC;
      xt_rsc_1_5_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_dp_inst_xt_rsc_1_5_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_dp_inst_xt_rsc_1_5_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_5_i_oswt => xt_rsc_1_5_i_oswt,
      xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_5_i_biwt => xt_rsc_1_5_i_biwt,
      xt_rsc_1_5_i_bdwt => xt_rsc_1_5_i_bdwt,
      xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_5_i_wea_d_core_sct_pff => xt_rsc_1_5_i_wea_d_core_sct_iff,
      xt_rsc_1_5_i_wea_d_core_psct_pff => xt_rsc_1_5_i_wea_d_core_psct_pff,
      xt_rsc_1_5_i_oswt_pff => xt_rsc_1_5_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_dp_inst : peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_5_i_qa_d => peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_dp_inst_xt_rsc_1_5_i_qa_d,
      xt_rsc_1_5_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_dp_inst_xt_rsc_1_5_i_qa_d_mxwt,
      xt_rsc_1_5_i_biwt => xt_rsc_1_5_i_biwt,
      xt_rsc_1_5_i_bdwt => xt_rsc_1_5_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_dp_inst_xt_rsc_1_5_i_qa_d <= xt_rsc_1_5_i_qa_d;
  xt_rsc_1_5_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_5_i_1_xt_rsc_1_5_wait_dp_inst_xt_rsc_1_5_i_qa_d_mxwt;

  xt_rsc_1_5_i_wea_d_pff <= xt_rsc_1_5_i_wea_d_core_sct_iff;
  xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_4_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_4_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_4_i_oswt : IN STD_LOGIC;
    xt_rsc_1_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_4_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_4_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_4_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_4_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_4_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_4_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_4_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_4_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_4_i_oswt : IN STD_LOGIC;
      xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_4_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_4_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_4_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_4_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_4_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_4_i_biwt : IN STD_LOGIC;
      xt_rsc_1_4_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_dp_inst_xt_rsc_1_4_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_dp_inst_xt_rsc_1_4_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_4_i_oswt => xt_rsc_1_4_i_oswt,
      xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_4_i_biwt => xt_rsc_1_4_i_biwt,
      xt_rsc_1_4_i_bdwt => xt_rsc_1_4_i_bdwt,
      xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_4_i_wea_d_core_sct_pff => xt_rsc_1_4_i_wea_d_core_sct_iff,
      xt_rsc_1_4_i_wea_d_core_psct_pff => xt_rsc_1_4_i_wea_d_core_psct_pff,
      xt_rsc_1_4_i_oswt_pff => xt_rsc_1_4_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_dp_inst : peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_4_i_qa_d => peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_dp_inst_xt_rsc_1_4_i_qa_d,
      xt_rsc_1_4_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_dp_inst_xt_rsc_1_4_i_qa_d_mxwt,
      xt_rsc_1_4_i_biwt => xt_rsc_1_4_i_biwt,
      xt_rsc_1_4_i_bdwt => xt_rsc_1_4_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_dp_inst_xt_rsc_1_4_i_qa_d <= xt_rsc_1_4_i_qa_d;
  xt_rsc_1_4_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_4_i_1_xt_rsc_1_4_wait_dp_inst_xt_rsc_1_4_i_qa_d_mxwt;

  xt_rsc_1_4_i_wea_d_pff <= xt_rsc_1_4_i_wea_d_core_sct_iff;
  xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_3_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_3_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_3_i_oswt : IN STD_LOGIC;
    xt_rsc_1_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_3_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_3_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_3_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_3_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_3_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_3_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_3_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_3_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_3_i_oswt : IN STD_LOGIC;
      xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_3_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_3_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_3_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_3_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_3_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_3_i_biwt : IN STD_LOGIC;
      xt_rsc_1_3_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_dp_inst_xt_rsc_1_3_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_dp_inst_xt_rsc_1_3_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_3_i_oswt => xt_rsc_1_3_i_oswt,
      xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_3_i_biwt => xt_rsc_1_3_i_biwt,
      xt_rsc_1_3_i_bdwt => xt_rsc_1_3_i_bdwt,
      xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_3_i_wea_d_core_sct_pff => xt_rsc_1_3_i_wea_d_core_sct_iff,
      xt_rsc_1_3_i_wea_d_core_psct_pff => xt_rsc_1_3_i_wea_d_core_psct_pff,
      xt_rsc_1_3_i_oswt_pff => xt_rsc_1_3_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_dp_inst : peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_3_i_qa_d => peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_dp_inst_xt_rsc_1_3_i_qa_d,
      xt_rsc_1_3_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_dp_inst_xt_rsc_1_3_i_qa_d_mxwt,
      xt_rsc_1_3_i_biwt => xt_rsc_1_3_i_biwt,
      xt_rsc_1_3_i_bdwt => xt_rsc_1_3_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_dp_inst_xt_rsc_1_3_i_qa_d <= xt_rsc_1_3_i_qa_d;
  xt_rsc_1_3_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_3_i_1_xt_rsc_1_3_wait_dp_inst_xt_rsc_1_3_i_qa_d_mxwt;

  xt_rsc_1_3_i_wea_d_pff <= xt_rsc_1_3_i_wea_d_core_sct_iff;
  xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_2_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_2_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_2_i_oswt : IN STD_LOGIC;
    xt_rsc_1_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_2_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_2_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_2_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_2_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_2_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_2_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_2_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_2_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_2_i_oswt : IN STD_LOGIC;
      xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_2_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_2_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_2_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_2_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_2_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_2_i_biwt : IN STD_LOGIC;
      xt_rsc_1_2_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_dp_inst_xt_rsc_1_2_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_dp_inst_xt_rsc_1_2_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_2_i_oswt => xt_rsc_1_2_i_oswt,
      xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_2_i_biwt => xt_rsc_1_2_i_biwt,
      xt_rsc_1_2_i_bdwt => xt_rsc_1_2_i_bdwt,
      xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_2_i_wea_d_core_sct_pff => xt_rsc_1_2_i_wea_d_core_sct_iff,
      xt_rsc_1_2_i_wea_d_core_psct_pff => xt_rsc_1_2_i_wea_d_core_psct_pff,
      xt_rsc_1_2_i_oswt_pff => xt_rsc_1_2_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_dp_inst : peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_2_i_qa_d => peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_dp_inst_xt_rsc_1_2_i_qa_d,
      xt_rsc_1_2_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_dp_inst_xt_rsc_1_2_i_qa_d_mxwt,
      xt_rsc_1_2_i_biwt => xt_rsc_1_2_i_biwt,
      xt_rsc_1_2_i_bdwt => xt_rsc_1_2_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_dp_inst_xt_rsc_1_2_i_qa_d <= xt_rsc_1_2_i_qa_d;
  xt_rsc_1_2_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_2_i_1_xt_rsc_1_2_wait_dp_inst_xt_rsc_1_2_i_qa_d_mxwt;

  xt_rsc_1_2_i_wea_d_pff <= xt_rsc_1_2_i_wea_d_core_sct_iff;
  xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_1_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_1_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_1_i_oswt : IN STD_LOGIC;
    xt_rsc_1_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_1_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_1_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_1_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_1_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_1_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_1_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_1_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_1_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_1_i_oswt : IN STD_LOGIC;
      xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_1_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_1_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_1_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_1_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_1_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_1_i_biwt : IN STD_LOGIC;
      xt_rsc_1_1_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_dp_inst_xt_rsc_1_1_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_dp_inst_xt_rsc_1_1_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_1_i_oswt => xt_rsc_1_1_i_oswt,
      xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_1_i_biwt => xt_rsc_1_1_i_biwt,
      xt_rsc_1_1_i_bdwt => xt_rsc_1_1_i_bdwt,
      xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_1_i_wea_d_core_sct_pff => xt_rsc_1_1_i_wea_d_core_sct_iff,
      xt_rsc_1_1_i_wea_d_core_psct_pff => xt_rsc_1_1_i_wea_d_core_psct_pff,
      xt_rsc_1_1_i_oswt_pff => xt_rsc_1_1_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_dp_inst : peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_1_i_qa_d => peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_dp_inst_xt_rsc_1_1_i_qa_d,
      xt_rsc_1_1_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_dp_inst_xt_rsc_1_1_i_qa_d_mxwt,
      xt_rsc_1_1_i_biwt => xt_rsc_1_1_i_biwt,
      xt_rsc_1_1_i_bdwt => xt_rsc_1_1_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_dp_inst_xt_rsc_1_1_i_qa_d <= xt_rsc_1_1_i_qa_d;
  xt_rsc_1_1_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_1_i_1_xt_rsc_1_1_wait_dp_inst_xt_rsc_1_1_i_qa_d_mxwt;

  xt_rsc_1_1_i_wea_d_pff <= xt_rsc_1_1_i_wea_d_core_sct_iff;
  xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_1_0_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_1_0_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_1_0_i_oswt : IN STD_LOGIC;
    xt_rsc_1_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_1_0_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_0_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_1_0_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_1_0_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_1_0_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_1_0_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_1_0_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_1_0_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_0_i_oswt : IN STD_LOGIC;
      xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_0_i_biwt : OUT STD_LOGIC;
      xt_rsc_1_0_i_bdwt : OUT STD_LOGIC;
      xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_1_0_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_1_0_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_0_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_0_i_biwt : IN STD_LOGIC;
      xt_rsc_1_0_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_dp_inst_xt_rsc_1_0_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_dp_inst_xt_rsc_1_0_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_ctrl_inst : peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_0_i_oswt => xt_rsc_1_0_i_oswt,
      xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_1_0_i_biwt => xt_rsc_1_0_i_biwt,
      xt_rsc_1_0_i_bdwt => xt_rsc_1_0_i_bdwt,
      xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_1_0_i_wea_d_core_sct_pff => xt_rsc_1_0_i_wea_d_core_sct_iff,
      xt_rsc_1_0_i_wea_d_core_psct_pff => xt_rsc_1_0_i_wea_d_core_psct_pff,
      xt_rsc_1_0_i_oswt_pff => xt_rsc_1_0_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_dp_inst : peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_0_i_qa_d => peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_dp_inst_xt_rsc_1_0_i_qa_d,
      xt_rsc_1_0_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_dp_inst_xt_rsc_1_0_i_qa_d_mxwt,
      xt_rsc_1_0_i_biwt => xt_rsc_1_0_i_biwt,
      xt_rsc_1_0_i_bdwt => xt_rsc_1_0_i_bdwt
    );
  peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_dp_inst_xt_rsc_1_0_i_qa_d <= xt_rsc_1_0_i_qa_d;
  xt_rsc_1_0_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_0_i_1_xt_rsc_1_0_wait_dp_inst_xt_rsc_1_0_i_qa_d_mxwt;

  xt_rsc_1_0_i_wea_d_pff <= xt_rsc_1_0_i_wea_d_core_sct_iff;
  xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_31_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_31_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_31_i_oswt : IN STD_LOGIC;
    xt_rsc_0_31_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_31_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_31_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_31_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_31_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_31_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_31_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_31_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_31_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_31_i_oswt : IN STD_LOGIC;
      xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_31_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_31_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_31_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_31_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_31_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_31_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_31_i_biwt : IN STD_LOGIC;
      xt_rsc_0_31_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_dp_inst_xt_rsc_0_31_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_dp_inst_xt_rsc_0_31_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_31_i_oswt => xt_rsc_0_31_i_oswt,
      xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_31_i_biwt => xt_rsc_0_31_i_biwt,
      xt_rsc_0_31_i_bdwt => xt_rsc_0_31_i_bdwt,
      xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_31_i_wea_d_core_sct_pff => xt_rsc_0_31_i_wea_d_core_sct_iff,
      xt_rsc_0_31_i_wea_d_core_psct_pff => xt_rsc_0_31_i_wea_d_core_psct_pff,
      xt_rsc_0_31_i_oswt_pff => xt_rsc_0_31_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_dp_inst : peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_31_i_qa_d => peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_dp_inst_xt_rsc_0_31_i_qa_d,
      xt_rsc_0_31_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_dp_inst_xt_rsc_0_31_i_qa_d_mxwt,
      xt_rsc_0_31_i_biwt => xt_rsc_0_31_i_biwt,
      xt_rsc_0_31_i_bdwt => xt_rsc_0_31_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_dp_inst_xt_rsc_0_31_i_qa_d <= xt_rsc_0_31_i_qa_d;
  xt_rsc_0_31_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_31_i_1_xt_rsc_0_31_wait_dp_inst_xt_rsc_0_31_i_qa_d_mxwt;

  xt_rsc_0_31_i_wea_d_pff <= xt_rsc_0_31_i_wea_d_core_sct_iff;
  xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_30_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_30_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_30_i_oswt : IN STD_LOGIC;
    xt_rsc_0_30_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_30_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_30_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_30_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_30_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_30_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_30_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_30_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_30_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_30_i_oswt : IN STD_LOGIC;
      xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_30_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_30_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_30_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_30_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_30_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_30_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_30_i_biwt : IN STD_LOGIC;
      xt_rsc_0_30_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_dp_inst_xt_rsc_0_30_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_dp_inst_xt_rsc_0_30_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_30_i_oswt => xt_rsc_0_30_i_oswt,
      xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_30_i_biwt => xt_rsc_0_30_i_biwt,
      xt_rsc_0_30_i_bdwt => xt_rsc_0_30_i_bdwt,
      xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_30_i_wea_d_core_sct_pff => xt_rsc_0_30_i_wea_d_core_sct_iff,
      xt_rsc_0_30_i_wea_d_core_psct_pff => xt_rsc_0_30_i_wea_d_core_psct_pff,
      xt_rsc_0_30_i_oswt_pff => xt_rsc_0_30_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_dp_inst : peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_30_i_qa_d => peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_dp_inst_xt_rsc_0_30_i_qa_d,
      xt_rsc_0_30_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_dp_inst_xt_rsc_0_30_i_qa_d_mxwt,
      xt_rsc_0_30_i_biwt => xt_rsc_0_30_i_biwt,
      xt_rsc_0_30_i_bdwt => xt_rsc_0_30_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_dp_inst_xt_rsc_0_30_i_qa_d <= xt_rsc_0_30_i_qa_d;
  xt_rsc_0_30_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_30_i_1_xt_rsc_0_30_wait_dp_inst_xt_rsc_0_30_i_qa_d_mxwt;

  xt_rsc_0_30_i_wea_d_pff <= xt_rsc_0_30_i_wea_d_core_sct_iff;
  xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_29_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_29_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_29_i_oswt : IN STD_LOGIC;
    xt_rsc_0_29_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_29_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_29_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_29_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_29_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_29_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_29_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_29_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_29_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_29_i_oswt : IN STD_LOGIC;
      xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_29_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_29_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_29_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_29_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_29_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_29_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_29_i_biwt : IN STD_LOGIC;
      xt_rsc_0_29_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_dp_inst_xt_rsc_0_29_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_dp_inst_xt_rsc_0_29_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_29_i_oswt => xt_rsc_0_29_i_oswt,
      xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_29_i_biwt => xt_rsc_0_29_i_biwt,
      xt_rsc_0_29_i_bdwt => xt_rsc_0_29_i_bdwt,
      xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_29_i_wea_d_core_sct_pff => xt_rsc_0_29_i_wea_d_core_sct_iff,
      xt_rsc_0_29_i_wea_d_core_psct_pff => xt_rsc_0_29_i_wea_d_core_psct_pff,
      xt_rsc_0_29_i_oswt_pff => xt_rsc_0_29_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_dp_inst : peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_29_i_qa_d => peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_dp_inst_xt_rsc_0_29_i_qa_d,
      xt_rsc_0_29_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_dp_inst_xt_rsc_0_29_i_qa_d_mxwt,
      xt_rsc_0_29_i_biwt => xt_rsc_0_29_i_biwt,
      xt_rsc_0_29_i_bdwt => xt_rsc_0_29_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_dp_inst_xt_rsc_0_29_i_qa_d <= xt_rsc_0_29_i_qa_d;
  xt_rsc_0_29_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_29_i_1_xt_rsc_0_29_wait_dp_inst_xt_rsc_0_29_i_qa_d_mxwt;

  xt_rsc_0_29_i_wea_d_pff <= xt_rsc_0_29_i_wea_d_core_sct_iff;
  xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_28_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_28_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_28_i_oswt : IN STD_LOGIC;
    xt_rsc_0_28_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_28_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_28_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_28_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_28_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_28_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_28_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_28_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_28_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_28_i_oswt : IN STD_LOGIC;
      xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_28_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_28_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_28_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_28_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_28_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_28_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_28_i_biwt : IN STD_LOGIC;
      xt_rsc_0_28_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_dp_inst_xt_rsc_0_28_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_dp_inst_xt_rsc_0_28_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_28_i_oswt => xt_rsc_0_28_i_oswt,
      xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_28_i_biwt => xt_rsc_0_28_i_biwt,
      xt_rsc_0_28_i_bdwt => xt_rsc_0_28_i_bdwt,
      xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_28_i_wea_d_core_sct_pff => xt_rsc_0_28_i_wea_d_core_sct_iff,
      xt_rsc_0_28_i_wea_d_core_psct_pff => xt_rsc_0_28_i_wea_d_core_psct_pff,
      xt_rsc_0_28_i_oswt_pff => xt_rsc_0_28_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_dp_inst : peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_28_i_qa_d => peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_dp_inst_xt_rsc_0_28_i_qa_d,
      xt_rsc_0_28_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_dp_inst_xt_rsc_0_28_i_qa_d_mxwt,
      xt_rsc_0_28_i_biwt => xt_rsc_0_28_i_biwt,
      xt_rsc_0_28_i_bdwt => xt_rsc_0_28_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_dp_inst_xt_rsc_0_28_i_qa_d <= xt_rsc_0_28_i_qa_d;
  xt_rsc_0_28_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_28_i_1_xt_rsc_0_28_wait_dp_inst_xt_rsc_0_28_i_qa_d_mxwt;

  xt_rsc_0_28_i_wea_d_pff <= xt_rsc_0_28_i_wea_d_core_sct_iff;
  xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_27_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_27_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_27_i_oswt : IN STD_LOGIC;
    xt_rsc_0_27_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_27_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_27_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_27_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_27_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_27_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_27_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_27_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_27_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_27_i_oswt : IN STD_LOGIC;
      xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_27_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_27_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_27_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_27_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_27_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_27_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_27_i_biwt : IN STD_LOGIC;
      xt_rsc_0_27_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_dp_inst_xt_rsc_0_27_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_dp_inst_xt_rsc_0_27_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_27_i_oswt => xt_rsc_0_27_i_oswt,
      xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_27_i_biwt => xt_rsc_0_27_i_biwt,
      xt_rsc_0_27_i_bdwt => xt_rsc_0_27_i_bdwt,
      xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_27_i_wea_d_core_sct_pff => xt_rsc_0_27_i_wea_d_core_sct_iff,
      xt_rsc_0_27_i_wea_d_core_psct_pff => xt_rsc_0_27_i_wea_d_core_psct_pff,
      xt_rsc_0_27_i_oswt_pff => xt_rsc_0_27_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_dp_inst : peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_27_i_qa_d => peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_dp_inst_xt_rsc_0_27_i_qa_d,
      xt_rsc_0_27_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_dp_inst_xt_rsc_0_27_i_qa_d_mxwt,
      xt_rsc_0_27_i_biwt => xt_rsc_0_27_i_biwt,
      xt_rsc_0_27_i_bdwt => xt_rsc_0_27_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_dp_inst_xt_rsc_0_27_i_qa_d <= xt_rsc_0_27_i_qa_d;
  xt_rsc_0_27_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_27_i_1_xt_rsc_0_27_wait_dp_inst_xt_rsc_0_27_i_qa_d_mxwt;

  xt_rsc_0_27_i_wea_d_pff <= xt_rsc_0_27_i_wea_d_core_sct_iff;
  xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_26_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_26_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_26_i_oswt : IN STD_LOGIC;
    xt_rsc_0_26_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_26_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_26_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_26_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_26_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_26_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_26_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_26_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_26_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_26_i_oswt : IN STD_LOGIC;
      xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_26_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_26_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_26_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_26_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_26_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_26_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_26_i_biwt : IN STD_LOGIC;
      xt_rsc_0_26_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_dp_inst_xt_rsc_0_26_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_dp_inst_xt_rsc_0_26_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_26_i_oswt => xt_rsc_0_26_i_oswt,
      xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_26_i_biwt => xt_rsc_0_26_i_biwt,
      xt_rsc_0_26_i_bdwt => xt_rsc_0_26_i_bdwt,
      xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_26_i_wea_d_core_sct_pff => xt_rsc_0_26_i_wea_d_core_sct_iff,
      xt_rsc_0_26_i_wea_d_core_psct_pff => xt_rsc_0_26_i_wea_d_core_psct_pff,
      xt_rsc_0_26_i_oswt_pff => xt_rsc_0_26_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_dp_inst : peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_26_i_qa_d => peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_dp_inst_xt_rsc_0_26_i_qa_d,
      xt_rsc_0_26_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_dp_inst_xt_rsc_0_26_i_qa_d_mxwt,
      xt_rsc_0_26_i_biwt => xt_rsc_0_26_i_biwt,
      xt_rsc_0_26_i_bdwt => xt_rsc_0_26_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_dp_inst_xt_rsc_0_26_i_qa_d <= xt_rsc_0_26_i_qa_d;
  xt_rsc_0_26_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_26_i_1_xt_rsc_0_26_wait_dp_inst_xt_rsc_0_26_i_qa_d_mxwt;

  xt_rsc_0_26_i_wea_d_pff <= xt_rsc_0_26_i_wea_d_core_sct_iff;
  xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_25_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_25_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_25_i_oswt : IN STD_LOGIC;
    xt_rsc_0_25_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_25_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_25_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_25_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_25_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_25_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_25_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_25_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_25_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_25_i_oswt : IN STD_LOGIC;
      xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_25_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_25_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_25_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_25_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_25_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_25_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_25_i_biwt : IN STD_LOGIC;
      xt_rsc_0_25_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_dp_inst_xt_rsc_0_25_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_dp_inst_xt_rsc_0_25_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_25_i_oswt => xt_rsc_0_25_i_oswt,
      xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_25_i_biwt => xt_rsc_0_25_i_biwt,
      xt_rsc_0_25_i_bdwt => xt_rsc_0_25_i_bdwt,
      xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_25_i_wea_d_core_sct_pff => xt_rsc_0_25_i_wea_d_core_sct_iff,
      xt_rsc_0_25_i_wea_d_core_psct_pff => xt_rsc_0_25_i_wea_d_core_psct_pff,
      xt_rsc_0_25_i_oswt_pff => xt_rsc_0_25_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_dp_inst : peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_25_i_qa_d => peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_dp_inst_xt_rsc_0_25_i_qa_d,
      xt_rsc_0_25_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_dp_inst_xt_rsc_0_25_i_qa_d_mxwt,
      xt_rsc_0_25_i_biwt => xt_rsc_0_25_i_biwt,
      xt_rsc_0_25_i_bdwt => xt_rsc_0_25_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_dp_inst_xt_rsc_0_25_i_qa_d <= xt_rsc_0_25_i_qa_d;
  xt_rsc_0_25_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_25_i_1_xt_rsc_0_25_wait_dp_inst_xt_rsc_0_25_i_qa_d_mxwt;

  xt_rsc_0_25_i_wea_d_pff <= xt_rsc_0_25_i_wea_d_core_sct_iff;
  xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_24_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_24_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_24_i_oswt : IN STD_LOGIC;
    xt_rsc_0_24_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_24_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_24_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_24_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_24_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_24_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_24_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_24_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_24_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_24_i_oswt : IN STD_LOGIC;
      xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_24_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_24_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_24_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_24_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_24_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_24_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_24_i_biwt : IN STD_LOGIC;
      xt_rsc_0_24_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_dp_inst_xt_rsc_0_24_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_dp_inst_xt_rsc_0_24_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_24_i_oswt => xt_rsc_0_24_i_oswt,
      xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_24_i_biwt => xt_rsc_0_24_i_biwt,
      xt_rsc_0_24_i_bdwt => xt_rsc_0_24_i_bdwt,
      xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_24_i_wea_d_core_sct_pff => xt_rsc_0_24_i_wea_d_core_sct_iff,
      xt_rsc_0_24_i_wea_d_core_psct_pff => xt_rsc_0_24_i_wea_d_core_psct_pff,
      xt_rsc_0_24_i_oswt_pff => xt_rsc_0_24_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_dp_inst : peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_24_i_qa_d => peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_dp_inst_xt_rsc_0_24_i_qa_d,
      xt_rsc_0_24_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_dp_inst_xt_rsc_0_24_i_qa_d_mxwt,
      xt_rsc_0_24_i_biwt => xt_rsc_0_24_i_biwt,
      xt_rsc_0_24_i_bdwt => xt_rsc_0_24_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_dp_inst_xt_rsc_0_24_i_qa_d <= xt_rsc_0_24_i_qa_d;
  xt_rsc_0_24_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_24_i_1_xt_rsc_0_24_wait_dp_inst_xt_rsc_0_24_i_qa_d_mxwt;

  xt_rsc_0_24_i_wea_d_pff <= xt_rsc_0_24_i_wea_d_core_sct_iff;
  xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_23_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_23_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_23_i_oswt : IN STD_LOGIC;
    xt_rsc_0_23_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_23_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_23_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_23_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_23_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_23_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_23_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_23_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_23_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_23_i_oswt : IN STD_LOGIC;
      xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_23_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_23_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_23_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_23_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_23_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_23_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_23_i_biwt : IN STD_LOGIC;
      xt_rsc_0_23_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_dp_inst_xt_rsc_0_23_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_dp_inst_xt_rsc_0_23_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_23_i_oswt => xt_rsc_0_23_i_oswt,
      xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_23_i_biwt => xt_rsc_0_23_i_biwt,
      xt_rsc_0_23_i_bdwt => xt_rsc_0_23_i_bdwt,
      xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_23_i_wea_d_core_sct_pff => xt_rsc_0_23_i_wea_d_core_sct_iff,
      xt_rsc_0_23_i_wea_d_core_psct_pff => xt_rsc_0_23_i_wea_d_core_psct_pff,
      xt_rsc_0_23_i_oswt_pff => xt_rsc_0_23_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_dp_inst : peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_23_i_qa_d => peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_dp_inst_xt_rsc_0_23_i_qa_d,
      xt_rsc_0_23_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_dp_inst_xt_rsc_0_23_i_qa_d_mxwt,
      xt_rsc_0_23_i_biwt => xt_rsc_0_23_i_biwt,
      xt_rsc_0_23_i_bdwt => xt_rsc_0_23_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_dp_inst_xt_rsc_0_23_i_qa_d <= xt_rsc_0_23_i_qa_d;
  xt_rsc_0_23_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_23_i_1_xt_rsc_0_23_wait_dp_inst_xt_rsc_0_23_i_qa_d_mxwt;

  xt_rsc_0_23_i_wea_d_pff <= xt_rsc_0_23_i_wea_d_core_sct_iff;
  xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_22_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_22_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_22_i_oswt : IN STD_LOGIC;
    xt_rsc_0_22_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_22_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_22_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_22_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_22_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_22_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_22_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_22_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_22_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_22_i_oswt : IN STD_LOGIC;
      xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_22_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_22_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_22_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_22_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_22_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_22_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_22_i_biwt : IN STD_LOGIC;
      xt_rsc_0_22_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_dp_inst_xt_rsc_0_22_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_dp_inst_xt_rsc_0_22_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_22_i_oswt => xt_rsc_0_22_i_oswt,
      xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_22_i_biwt => xt_rsc_0_22_i_biwt,
      xt_rsc_0_22_i_bdwt => xt_rsc_0_22_i_bdwt,
      xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_22_i_wea_d_core_sct_pff => xt_rsc_0_22_i_wea_d_core_sct_iff,
      xt_rsc_0_22_i_wea_d_core_psct_pff => xt_rsc_0_22_i_wea_d_core_psct_pff,
      xt_rsc_0_22_i_oswt_pff => xt_rsc_0_22_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_dp_inst : peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_22_i_qa_d => peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_dp_inst_xt_rsc_0_22_i_qa_d,
      xt_rsc_0_22_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_dp_inst_xt_rsc_0_22_i_qa_d_mxwt,
      xt_rsc_0_22_i_biwt => xt_rsc_0_22_i_biwt,
      xt_rsc_0_22_i_bdwt => xt_rsc_0_22_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_dp_inst_xt_rsc_0_22_i_qa_d <= xt_rsc_0_22_i_qa_d;
  xt_rsc_0_22_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_22_i_1_xt_rsc_0_22_wait_dp_inst_xt_rsc_0_22_i_qa_d_mxwt;

  xt_rsc_0_22_i_wea_d_pff <= xt_rsc_0_22_i_wea_d_core_sct_iff;
  xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_21_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_21_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_21_i_oswt : IN STD_LOGIC;
    xt_rsc_0_21_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_21_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_21_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_21_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_21_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_21_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_21_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_21_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_21_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_21_i_oswt : IN STD_LOGIC;
      xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_21_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_21_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_21_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_21_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_21_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_21_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_21_i_biwt : IN STD_LOGIC;
      xt_rsc_0_21_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_dp_inst_xt_rsc_0_21_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_dp_inst_xt_rsc_0_21_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_21_i_oswt => xt_rsc_0_21_i_oswt,
      xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_21_i_biwt => xt_rsc_0_21_i_biwt,
      xt_rsc_0_21_i_bdwt => xt_rsc_0_21_i_bdwt,
      xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_21_i_wea_d_core_sct_pff => xt_rsc_0_21_i_wea_d_core_sct_iff,
      xt_rsc_0_21_i_wea_d_core_psct_pff => xt_rsc_0_21_i_wea_d_core_psct_pff,
      xt_rsc_0_21_i_oswt_pff => xt_rsc_0_21_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_dp_inst : peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_21_i_qa_d => peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_dp_inst_xt_rsc_0_21_i_qa_d,
      xt_rsc_0_21_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_dp_inst_xt_rsc_0_21_i_qa_d_mxwt,
      xt_rsc_0_21_i_biwt => xt_rsc_0_21_i_biwt,
      xt_rsc_0_21_i_bdwt => xt_rsc_0_21_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_dp_inst_xt_rsc_0_21_i_qa_d <= xt_rsc_0_21_i_qa_d;
  xt_rsc_0_21_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_21_i_1_xt_rsc_0_21_wait_dp_inst_xt_rsc_0_21_i_qa_d_mxwt;

  xt_rsc_0_21_i_wea_d_pff <= xt_rsc_0_21_i_wea_d_core_sct_iff;
  xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_20_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_20_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_20_i_oswt : IN STD_LOGIC;
    xt_rsc_0_20_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_20_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_20_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_20_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_20_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_20_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_20_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_20_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_20_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_20_i_oswt : IN STD_LOGIC;
      xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_20_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_20_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_20_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_20_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_20_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_20_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_20_i_biwt : IN STD_LOGIC;
      xt_rsc_0_20_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_dp_inst_xt_rsc_0_20_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_dp_inst_xt_rsc_0_20_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_20_i_oswt => xt_rsc_0_20_i_oswt,
      xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_20_i_biwt => xt_rsc_0_20_i_biwt,
      xt_rsc_0_20_i_bdwt => xt_rsc_0_20_i_bdwt,
      xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_20_i_wea_d_core_sct_pff => xt_rsc_0_20_i_wea_d_core_sct_iff,
      xt_rsc_0_20_i_wea_d_core_psct_pff => xt_rsc_0_20_i_wea_d_core_psct_pff,
      xt_rsc_0_20_i_oswt_pff => xt_rsc_0_20_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_dp_inst : peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_20_i_qa_d => peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_dp_inst_xt_rsc_0_20_i_qa_d,
      xt_rsc_0_20_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_dp_inst_xt_rsc_0_20_i_qa_d_mxwt,
      xt_rsc_0_20_i_biwt => xt_rsc_0_20_i_biwt,
      xt_rsc_0_20_i_bdwt => xt_rsc_0_20_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_dp_inst_xt_rsc_0_20_i_qa_d <= xt_rsc_0_20_i_qa_d;
  xt_rsc_0_20_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_20_i_1_xt_rsc_0_20_wait_dp_inst_xt_rsc_0_20_i_qa_d_mxwt;

  xt_rsc_0_20_i_wea_d_pff <= xt_rsc_0_20_i_wea_d_core_sct_iff;
  xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_19_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_19_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_19_i_oswt : IN STD_LOGIC;
    xt_rsc_0_19_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_19_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_19_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_19_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_19_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_19_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_19_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_19_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_19_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_19_i_oswt : IN STD_LOGIC;
      xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_19_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_19_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_19_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_19_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_19_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_19_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_19_i_biwt : IN STD_LOGIC;
      xt_rsc_0_19_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_dp_inst_xt_rsc_0_19_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_dp_inst_xt_rsc_0_19_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_19_i_oswt => xt_rsc_0_19_i_oswt,
      xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_19_i_biwt => xt_rsc_0_19_i_biwt,
      xt_rsc_0_19_i_bdwt => xt_rsc_0_19_i_bdwt,
      xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_19_i_wea_d_core_sct_pff => xt_rsc_0_19_i_wea_d_core_sct_iff,
      xt_rsc_0_19_i_wea_d_core_psct_pff => xt_rsc_0_19_i_wea_d_core_psct_pff,
      xt_rsc_0_19_i_oswt_pff => xt_rsc_0_19_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_dp_inst : peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_19_i_qa_d => peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_dp_inst_xt_rsc_0_19_i_qa_d,
      xt_rsc_0_19_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_dp_inst_xt_rsc_0_19_i_qa_d_mxwt,
      xt_rsc_0_19_i_biwt => xt_rsc_0_19_i_biwt,
      xt_rsc_0_19_i_bdwt => xt_rsc_0_19_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_dp_inst_xt_rsc_0_19_i_qa_d <= xt_rsc_0_19_i_qa_d;
  xt_rsc_0_19_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_19_i_1_xt_rsc_0_19_wait_dp_inst_xt_rsc_0_19_i_qa_d_mxwt;

  xt_rsc_0_19_i_wea_d_pff <= xt_rsc_0_19_i_wea_d_core_sct_iff;
  xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_18_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_18_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_18_i_oswt : IN STD_LOGIC;
    xt_rsc_0_18_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_18_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_18_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_18_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_18_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_18_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_18_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_18_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_18_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_18_i_oswt : IN STD_LOGIC;
      xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_18_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_18_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_18_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_18_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_18_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_18_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_18_i_biwt : IN STD_LOGIC;
      xt_rsc_0_18_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_dp_inst_xt_rsc_0_18_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_dp_inst_xt_rsc_0_18_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_18_i_oswt => xt_rsc_0_18_i_oswt,
      xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_18_i_biwt => xt_rsc_0_18_i_biwt,
      xt_rsc_0_18_i_bdwt => xt_rsc_0_18_i_bdwt,
      xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_18_i_wea_d_core_sct_pff => xt_rsc_0_18_i_wea_d_core_sct_iff,
      xt_rsc_0_18_i_wea_d_core_psct_pff => xt_rsc_0_18_i_wea_d_core_psct_pff,
      xt_rsc_0_18_i_oswt_pff => xt_rsc_0_18_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_dp_inst : peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_18_i_qa_d => peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_dp_inst_xt_rsc_0_18_i_qa_d,
      xt_rsc_0_18_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_dp_inst_xt_rsc_0_18_i_qa_d_mxwt,
      xt_rsc_0_18_i_biwt => xt_rsc_0_18_i_biwt,
      xt_rsc_0_18_i_bdwt => xt_rsc_0_18_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_dp_inst_xt_rsc_0_18_i_qa_d <= xt_rsc_0_18_i_qa_d;
  xt_rsc_0_18_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_18_i_1_xt_rsc_0_18_wait_dp_inst_xt_rsc_0_18_i_qa_d_mxwt;

  xt_rsc_0_18_i_wea_d_pff <= xt_rsc_0_18_i_wea_d_core_sct_iff;
  xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_17_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_17_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_17_i_oswt : IN STD_LOGIC;
    xt_rsc_0_17_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_17_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_17_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_17_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_17_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_17_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_17_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_17_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_17_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_17_i_oswt : IN STD_LOGIC;
      xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_17_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_17_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_17_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_17_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_17_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_17_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_17_i_biwt : IN STD_LOGIC;
      xt_rsc_0_17_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_dp_inst_xt_rsc_0_17_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_dp_inst_xt_rsc_0_17_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_17_i_oswt => xt_rsc_0_17_i_oswt,
      xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_17_i_biwt => xt_rsc_0_17_i_biwt,
      xt_rsc_0_17_i_bdwt => xt_rsc_0_17_i_bdwt,
      xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_17_i_wea_d_core_sct_pff => xt_rsc_0_17_i_wea_d_core_sct_iff,
      xt_rsc_0_17_i_wea_d_core_psct_pff => xt_rsc_0_17_i_wea_d_core_psct_pff,
      xt_rsc_0_17_i_oswt_pff => xt_rsc_0_17_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_dp_inst : peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_17_i_qa_d => peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_dp_inst_xt_rsc_0_17_i_qa_d,
      xt_rsc_0_17_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_dp_inst_xt_rsc_0_17_i_qa_d_mxwt,
      xt_rsc_0_17_i_biwt => xt_rsc_0_17_i_biwt,
      xt_rsc_0_17_i_bdwt => xt_rsc_0_17_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_dp_inst_xt_rsc_0_17_i_qa_d <= xt_rsc_0_17_i_qa_d;
  xt_rsc_0_17_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_17_i_1_xt_rsc_0_17_wait_dp_inst_xt_rsc_0_17_i_qa_d_mxwt;

  xt_rsc_0_17_i_wea_d_pff <= xt_rsc_0_17_i_wea_d_core_sct_iff;
  xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_16_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_16_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_16_i_oswt : IN STD_LOGIC;
    xt_rsc_0_16_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_16_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_16_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_16_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_16_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_16_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_16_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_16_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_16_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_16_i_oswt : IN STD_LOGIC;
      xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_16_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_16_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_16_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_16_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_16_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_16_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_16_i_biwt : IN STD_LOGIC;
      xt_rsc_0_16_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_dp_inst_xt_rsc_0_16_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_dp_inst_xt_rsc_0_16_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_16_i_oswt => xt_rsc_0_16_i_oswt,
      xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_16_i_biwt => xt_rsc_0_16_i_biwt,
      xt_rsc_0_16_i_bdwt => xt_rsc_0_16_i_bdwt,
      xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_16_i_wea_d_core_sct_pff => xt_rsc_0_16_i_wea_d_core_sct_iff,
      xt_rsc_0_16_i_wea_d_core_psct_pff => xt_rsc_0_16_i_wea_d_core_psct_pff,
      xt_rsc_0_16_i_oswt_pff => xt_rsc_0_16_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_dp_inst : peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_16_i_qa_d => peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_dp_inst_xt_rsc_0_16_i_qa_d,
      xt_rsc_0_16_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_dp_inst_xt_rsc_0_16_i_qa_d_mxwt,
      xt_rsc_0_16_i_biwt => xt_rsc_0_16_i_biwt,
      xt_rsc_0_16_i_bdwt => xt_rsc_0_16_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_dp_inst_xt_rsc_0_16_i_qa_d <= xt_rsc_0_16_i_qa_d;
  xt_rsc_0_16_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_16_i_1_xt_rsc_0_16_wait_dp_inst_xt_rsc_0_16_i_qa_d_mxwt;

  xt_rsc_0_16_i_wea_d_pff <= xt_rsc_0_16_i_wea_d_core_sct_iff;
  xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_15_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_15_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_15_i_oswt : IN STD_LOGIC;
    xt_rsc_0_15_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_15_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_15_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_15_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_15_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_15_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_15_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_15_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_15_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_15_i_oswt : IN STD_LOGIC;
      xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_15_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_15_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_15_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_15_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_15_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_15_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_15_i_biwt : IN STD_LOGIC;
      xt_rsc_0_15_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_dp_inst_xt_rsc_0_15_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_dp_inst_xt_rsc_0_15_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_15_i_oswt => xt_rsc_0_15_i_oswt,
      xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_15_i_biwt => xt_rsc_0_15_i_biwt,
      xt_rsc_0_15_i_bdwt => xt_rsc_0_15_i_bdwt,
      xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_15_i_wea_d_core_sct_pff => xt_rsc_0_15_i_wea_d_core_sct_iff,
      xt_rsc_0_15_i_wea_d_core_psct_pff => xt_rsc_0_15_i_wea_d_core_psct_pff,
      xt_rsc_0_15_i_oswt_pff => xt_rsc_0_15_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_dp_inst : peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_15_i_qa_d => peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_dp_inst_xt_rsc_0_15_i_qa_d,
      xt_rsc_0_15_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_dp_inst_xt_rsc_0_15_i_qa_d_mxwt,
      xt_rsc_0_15_i_biwt => xt_rsc_0_15_i_biwt,
      xt_rsc_0_15_i_bdwt => xt_rsc_0_15_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_dp_inst_xt_rsc_0_15_i_qa_d <= xt_rsc_0_15_i_qa_d;
  xt_rsc_0_15_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_15_i_1_xt_rsc_0_15_wait_dp_inst_xt_rsc_0_15_i_qa_d_mxwt;

  xt_rsc_0_15_i_wea_d_pff <= xt_rsc_0_15_i_wea_d_core_sct_iff;
  xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_14_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_14_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_14_i_oswt : IN STD_LOGIC;
    xt_rsc_0_14_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_14_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_14_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_14_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_14_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_14_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_14_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_14_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_14_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_14_i_oswt : IN STD_LOGIC;
      xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_14_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_14_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_14_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_14_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_14_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_14_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_14_i_biwt : IN STD_LOGIC;
      xt_rsc_0_14_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_dp_inst_xt_rsc_0_14_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_dp_inst_xt_rsc_0_14_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_14_i_oswt => xt_rsc_0_14_i_oswt,
      xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_14_i_biwt => xt_rsc_0_14_i_biwt,
      xt_rsc_0_14_i_bdwt => xt_rsc_0_14_i_bdwt,
      xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_14_i_wea_d_core_sct_pff => xt_rsc_0_14_i_wea_d_core_sct_iff,
      xt_rsc_0_14_i_wea_d_core_psct_pff => xt_rsc_0_14_i_wea_d_core_psct_pff,
      xt_rsc_0_14_i_oswt_pff => xt_rsc_0_14_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_dp_inst : peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_14_i_qa_d => peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_dp_inst_xt_rsc_0_14_i_qa_d,
      xt_rsc_0_14_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_dp_inst_xt_rsc_0_14_i_qa_d_mxwt,
      xt_rsc_0_14_i_biwt => xt_rsc_0_14_i_biwt,
      xt_rsc_0_14_i_bdwt => xt_rsc_0_14_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_dp_inst_xt_rsc_0_14_i_qa_d <= xt_rsc_0_14_i_qa_d;
  xt_rsc_0_14_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_14_i_1_xt_rsc_0_14_wait_dp_inst_xt_rsc_0_14_i_qa_d_mxwt;

  xt_rsc_0_14_i_wea_d_pff <= xt_rsc_0_14_i_wea_d_core_sct_iff;
  xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_13_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_13_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_13_i_oswt : IN STD_LOGIC;
    xt_rsc_0_13_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_13_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_13_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_13_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_13_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_13_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_13_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_13_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_13_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_13_i_oswt : IN STD_LOGIC;
      xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_13_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_13_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_13_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_13_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_13_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_13_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_13_i_biwt : IN STD_LOGIC;
      xt_rsc_0_13_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_dp_inst_xt_rsc_0_13_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_dp_inst_xt_rsc_0_13_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_13_i_oswt => xt_rsc_0_13_i_oswt,
      xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_13_i_biwt => xt_rsc_0_13_i_biwt,
      xt_rsc_0_13_i_bdwt => xt_rsc_0_13_i_bdwt,
      xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_13_i_wea_d_core_sct_pff => xt_rsc_0_13_i_wea_d_core_sct_iff,
      xt_rsc_0_13_i_wea_d_core_psct_pff => xt_rsc_0_13_i_wea_d_core_psct_pff,
      xt_rsc_0_13_i_oswt_pff => xt_rsc_0_13_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_dp_inst : peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_13_i_qa_d => peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_dp_inst_xt_rsc_0_13_i_qa_d,
      xt_rsc_0_13_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_dp_inst_xt_rsc_0_13_i_qa_d_mxwt,
      xt_rsc_0_13_i_biwt => xt_rsc_0_13_i_biwt,
      xt_rsc_0_13_i_bdwt => xt_rsc_0_13_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_dp_inst_xt_rsc_0_13_i_qa_d <= xt_rsc_0_13_i_qa_d;
  xt_rsc_0_13_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_13_i_1_xt_rsc_0_13_wait_dp_inst_xt_rsc_0_13_i_qa_d_mxwt;

  xt_rsc_0_13_i_wea_d_pff <= xt_rsc_0_13_i_wea_d_core_sct_iff;
  xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_12_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_12_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_12_i_oswt : IN STD_LOGIC;
    xt_rsc_0_12_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_12_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_12_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_12_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_12_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_12_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_12_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_12_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_12_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_12_i_oswt : IN STD_LOGIC;
      xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_12_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_12_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_12_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_12_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_12_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_12_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_12_i_biwt : IN STD_LOGIC;
      xt_rsc_0_12_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_dp_inst_xt_rsc_0_12_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_dp_inst_xt_rsc_0_12_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_12_i_oswt => xt_rsc_0_12_i_oswt,
      xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_12_i_biwt => xt_rsc_0_12_i_biwt,
      xt_rsc_0_12_i_bdwt => xt_rsc_0_12_i_bdwt,
      xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_12_i_wea_d_core_sct_pff => xt_rsc_0_12_i_wea_d_core_sct_iff,
      xt_rsc_0_12_i_wea_d_core_psct_pff => xt_rsc_0_12_i_wea_d_core_psct_pff,
      xt_rsc_0_12_i_oswt_pff => xt_rsc_0_12_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_dp_inst : peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_12_i_qa_d => peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_dp_inst_xt_rsc_0_12_i_qa_d,
      xt_rsc_0_12_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_dp_inst_xt_rsc_0_12_i_qa_d_mxwt,
      xt_rsc_0_12_i_biwt => xt_rsc_0_12_i_biwt,
      xt_rsc_0_12_i_bdwt => xt_rsc_0_12_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_dp_inst_xt_rsc_0_12_i_qa_d <= xt_rsc_0_12_i_qa_d;
  xt_rsc_0_12_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_12_i_1_xt_rsc_0_12_wait_dp_inst_xt_rsc_0_12_i_qa_d_mxwt;

  xt_rsc_0_12_i_wea_d_pff <= xt_rsc_0_12_i_wea_d_core_sct_iff;
  xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_11_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_11_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_11_i_oswt : IN STD_LOGIC;
    xt_rsc_0_11_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_11_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_11_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_11_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_11_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_11_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_11_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_11_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_11_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_11_i_oswt : IN STD_LOGIC;
      xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_11_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_11_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_11_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_11_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_11_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_11_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_11_i_biwt : IN STD_LOGIC;
      xt_rsc_0_11_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_dp_inst_xt_rsc_0_11_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_dp_inst_xt_rsc_0_11_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_11_i_oswt => xt_rsc_0_11_i_oswt,
      xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_11_i_biwt => xt_rsc_0_11_i_biwt,
      xt_rsc_0_11_i_bdwt => xt_rsc_0_11_i_bdwt,
      xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_11_i_wea_d_core_sct_pff => xt_rsc_0_11_i_wea_d_core_sct_iff,
      xt_rsc_0_11_i_wea_d_core_psct_pff => xt_rsc_0_11_i_wea_d_core_psct_pff,
      xt_rsc_0_11_i_oswt_pff => xt_rsc_0_11_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_dp_inst : peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_11_i_qa_d => peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_dp_inst_xt_rsc_0_11_i_qa_d,
      xt_rsc_0_11_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_dp_inst_xt_rsc_0_11_i_qa_d_mxwt,
      xt_rsc_0_11_i_biwt => xt_rsc_0_11_i_biwt,
      xt_rsc_0_11_i_bdwt => xt_rsc_0_11_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_dp_inst_xt_rsc_0_11_i_qa_d <= xt_rsc_0_11_i_qa_d;
  xt_rsc_0_11_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_11_i_1_xt_rsc_0_11_wait_dp_inst_xt_rsc_0_11_i_qa_d_mxwt;

  xt_rsc_0_11_i_wea_d_pff <= xt_rsc_0_11_i_wea_d_core_sct_iff;
  xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_10_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_10_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_10_i_oswt : IN STD_LOGIC;
    xt_rsc_0_10_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_10_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_10_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_10_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_10_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_10_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_10_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_10_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_10_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_10_i_oswt : IN STD_LOGIC;
      xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_10_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_10_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_10_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_10_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_10_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_10_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_10_i_biwt : IN STD_LOGIC;
      xt_rsc_0_10_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_dp_inst_xt_rsc_0_10_i_qa_d
      : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_dp_inst_xt_rsc_0_10_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_10_i_oswt => xt_rsc_0_10_i_oswt,
      xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_10_i_biwt => xt_rsc_0_10_i_biwt,
      xt_rsc_0_10_i_bdwt => xt_rsc_0_10_i_bdwt,
      xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_10_i_wea_d_core_sct_pff => xt_rsc_0_10_i_wea_d_core_sct_iff,
      xt_rsc_0_10_i_wea_d_core_psct_pff => xt_rsc_0_10_i_wea_d_core_psct_pff,
      xt_rsc_0_10_i_oswt_pff => xt_rsc_0_10_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_dp_inst : peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_10_i_qa_d => peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_dp_inst_xt_rsc_0_10_i_qa_d,
      xt_rsc_0_10_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_dp_inst_xt_rsc_0_10_i_qa_d_mxwt,
      xt_rsc_0_10_i_biwt => xt_rsc_0_10_i_biwt,
      xt_rsc_0_10_i_bdwt => xt_rsc_0_10_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_dp_inst_xt_rsc_0_10_i_qa_d <= xt_rsc_0_10_i_qa_d;
  xt_rsc_0_10_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_10_i_1_xt_rsc_0_10_wait_dp_inst_xt_rsc_0_10_i_qa_d_mxwt;

  xt_rsc_0_10_i_wea_d_pff <= xt_rsc_0_10_i_wea_d_core_sct_iff;
  xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_9_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_9_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_9_i_oswt : IN STD_LOGIC;
    xt_rsc_0_9_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_9_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_9_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_9_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_9_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_9_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_9_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_9_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_9_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_9_i_oswt : IN STD_LOGIC;
      xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_9_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_9_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_9_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_9_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_9_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_9_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_9_i_biwt : IN STD_LOGIC;
      xt_rsc_0_9_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_dp_inst_xt_rsc_0_9_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_dp_inst_xt_rsc_0_9_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_9_i_oswt => xt_rsc_0_9_i_oswt,
      xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_9_i_biwt => xt_rsc_0_9_i_biwt,
      xt_rsc_0_9_i_bdwt => xt_rsc_0_9_i_bdwt,
      xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_9_i_wea_d_core_sct_pff => xt_rsc_0_9_i_wea_d_core_sct_iff,
      xt_rsc_0_9_i_wea_d_core_psct_pff => xt_rsc_0_9_i_wea_d_core_psct_pff,
      xt_rsc_0_9_i_oswt_pff => xt_rsc_0_9_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_dp_inst : peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_9_i_qa_d => peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_dp_inst_xt_rsc_0_9_i_qa_d,
      xt_rsc_0_9_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_dp_inst_xt_rsc_0_9_i_qa_d_mxwt,
      xt_rsc_0_9_i_biwt => xt_rsc_0_9_i_biwt,
      xt_rsc_0_9_i_bdwt => xt_rsc_0_9_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_dp_inst_xt_rsc_0_9_i_qa_d <= xt_rsc_0_9_i_qa_d;
  xt_rsc_0_9_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_9_i_1_xt_rsc_0_9_wait_dp_inst_xt_rsc_0_9_i_qa_d_mxwt;

  xt_rsc_0_9_i_wea_d_pff <= xt_rsc_0_9_i_wea_d_core_sct_iff;
  xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_8_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_8_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_8_i_oswt : IN STD_LOGIC;
    xt_rsc_0_8_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_8_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_8_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_8_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_8_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_8_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_8_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_8_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_8_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_8_i_oswt : IN STD_LOGIC;
      xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_8_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_8_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_8_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_8_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_8_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_8_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_8_i_biwt : IN STD_LOGIC;
      xt_rsc_0_8_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_dp_inst_xt_rsc_0_8_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_dp_inst_xt_rsc_0_8_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_8_i_oswt => xt_rsc_0_8_i_oswt,
      xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_8_i_biwt => xt_rsc_0_8_i_biwt,
      xt_rsc_0_8_i_bdwt => xt_rsc_0_8_i_bdwt,
      xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_8_i_wea_d_core_sct_pff => xt_rsc_0_8_i_wea_d_core_sct_iff,
      xt_rsc_0_8_i_wea_d_core_psct_pff => xt_rsc_0_8_i_wea_d_core_psct_pff,
      xt_rsc_0_8_i_oswt_pff => xt_rsc_0_8_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_dp_inst : peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_8_i_qa_d => peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_dp_inst_xt_rsc_0_8_i_qa_d,
      xt_rsc_0_8_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_dp_inst_xt_rsc_0_8_i_qa_d_mxwt,
      xt_rsc_0_8_i_biwt => xt_rsc_0_8_i_biwt,
      xt_rsc_0_8_i_bdwt => xt_rsc_0_8_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_dp_inst_xt_rsc_0_8_i_qa_d <= xt_rsc_0_8_i_qa_d;
  xt_rsc_0_8_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_8_i_1_xt_rsc_0_8_wait_dp_inst_xt_rsc_0_8_i_qa_d_mxwt;

  xt_rsc_0_8_i_wea_d_pff <= xt_rsc_0_8_i_wea_d_core_sct_iff;
  xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_7_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_7_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_7_i_oswt : IN STD_LOGIC;
    xt_rsc_0_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_7_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_7_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_7_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_7_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_7_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_7_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_7_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_7_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_7_i_oswt : IN STD_LOGIC;
      xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_7_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_7_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_7_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_7_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_7_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_7_i_biwt : IN STD_LOGIC;
      xt_rsc_0_7_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_dp_inst_xt_rsc_0_7_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_dp_inst_xt_rsc_0_7_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_7_i_oswt => xt_rsc_0_7_i_oswt,
      xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_7_i_biwt => xt_rsc_0_7_i_biwt,
      xt_rsc_0_7_i_bdwt => xt_rsc_0_7_i_bdwt,
      xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_7_i_wea_d_core_sct_pff => xt_rsc_0_7_i_wea_d_core_sct_iff,
      xt_rsc_0_7_i_wea_d_core_psct_pff => xt_rsc_0_7_i_wea_d_core_psct_pff,
      xt_rsc_0_7_i_oswt_pff => xt_rsc_0_7_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_dp_inst : peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_7_i_qa_d => peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_dp_inst_xt_rsc_0_7_i_qa_d,
      xt_rsc_0_7_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_dp_inst_xt_rsc_0_7_i_qa_d_mxwt,
      xt_rsc_0_7_i_biwt => xt_rsc_0_7_i_biwt,
      xt_rsc_0_7_i_bdwt => xt_rsc_0_7_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_dp_inst_xt_rsc_0_7_i_qa_d <= xt_rsc_0_7_i_qa_d;
  xt_rsc_0_7_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_7_i_1_xt_rsc_0_7_wait_dp_inst_xt_rsc_0_7_i_qa_d_mxwt;

  xt_rsc_0_7_i_wea_d_pff <= xt_rsc_0_7_i_wea_d_core_sct_iff;
  xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_6_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_6_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_6_i_oswt : IN STD_LOGIC;
    xt_rsc_0_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_6_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_6_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_6_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_6_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_6_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_6_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_6_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_6_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_6_i_oswt : IN STD_LOGIC;
      xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_6_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_6_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_6_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_6_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_6_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_6_i_biwt : IN STD_LOGIC;
      xt_rsc_0_6_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_dp_inst_xt_rsc_0_6_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_dp_inst_xt_rsc_0_6_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_6_i_oswt => xt_rsc_0_6_i_oswt,
      xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_6_i_biwt => xt_rsc_0_6_i_biwt,
      xt_rsc_0_6_i_bdwt => xt_rsc_0_6_i_bdwt,
      xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_6_i_wea_d_core_sct_pff => xt_rsc_0_6_i_wea_d_core_sct_iff,
      xt_rsc_0_6_i_wea_d_core_psct_pff => xt_rsc_0_6_i_wea_d_core_psct_pff,
      xt_rsc_0_6_i_oswt_pff => xt_rsc_0_6_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_dp_inst : peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_6_i_qa_d => peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_dp_inst_xt_rsc_0_6_i_qa_d,
      xt_rsc_0_6_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_dp_inst_xt_rsc_0_6_i_qa_d_mxwt,
      xt_rsc_0_6_i_biwt => xt_rsc_0_6_i_biwt,
      xt_rsc_0_6_i_bdwt => xt_rsc_0_6_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_dp_inst_xt_rsc_0_6_i_qa_d <= xt_rsc_0_6_i_qa_d;
  xt_rsc_0_6_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_6_i_1_xt_rsc_0_6_wait_dp_inst_xt_rsc_0_6_i_qa_d_mxwt;

  xt_rsc_0_6_i_wea_d_pff <= xt_rsc_0_6_i_wea_d_core_sct_iff;
  xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_5_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_5_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_5_i_oswt : IN STD_LOGIC;
    xt_rsc_0_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_5_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_5_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_5_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_5_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_5_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_5_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_5_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_5_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_5_i_oswt : IN STD_LOGIC;
      xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_5_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_5_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_5_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_5_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_5_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_5_i_biwt : IN STD_LOGIC;
      xt_rsc_0_5_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_dp_inst_xt_rsc_0_5_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_dp_inst_xt_rsc_0_5_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_5_i_oswt => xt_rsc_0_5_i_oswt,
      xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_5_i_biwt => xt_rsc_0_5_i_biwt,
      xt_rsc_0_5_i_bdwt => xt_rsc_0_5_i_bdwt,
      xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_5_i_wea_d_core_sct_pff => xt_rsc_0_5_i_wea_d_core_sct_iff,
      xt_rsc_0_5_i_wea_d_core_psct_pff => xt_rsc_0_5_i_wea_d_core_psct_pff,
      xt_rsc_0_5_i_oswt_pff => xt_rsc_0_5_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_dp_inst : peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_5_i_qa_d => peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_dp_inst_xt_rsc_0_5_i_qa_d,
      xt_rsc_0_5_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_dp_inst_xt_rsc_0_5_i_qa_d_mxwt,
      xt_rsc_0_5_i_biwt => xt_rsc_0_5_i_biwt,
      xt_rsc_0_5_i_bdwt => xt_rsc_0_5_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_dp_inst_xt_rsc_0_5_i_qa_d <= xt_rsc_0_5_i_qa_d;
  xt_rsc_0_5_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_5_i_1_xt_rsc_0_5_wait_dp_inst_xt_rsc_0_5_i_qa_d_mxwt;

  xt_rsc_0_5_i_wea_d_pff <= xt_rsc_0_5_i_wea_d_core_sct_iff;
  xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_4_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_4_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_4_i_oswt : IN STD_LOGIC;
    xt_rsc_0_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_4_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_4_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_4_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_4_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_4_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_4_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_4_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_4_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_4_i_oswt : IN STD_LOGIC;
      xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_4_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_4_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_4_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_4_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_4_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_4_i_biwt : IN STD_LOGIC;
      xt_rsc_0_4_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_dp_inst_xt_rsc_0_4_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_dp_inst_xt_rsc_0_4_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_4_i_oswt => xt_rsc_0_4_i_oswt,
      xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_4_i_biwt => xt_rsc_0_4_i_biwt,
      xt_rsc_0_4_i_bdwt => xt_rsc_0_4_i_bdwt,
      xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_4_i_wea_d_core_sct_pff => xt_rsc_0_4_i_wea_d_core_sct_iff,
      xt_rsc_0_4_i_wea_d_core_psct_pff => xt_rsc_0_4_i_wea_d_core_psct_pff,
      xt_rsc_0_4_i_oswt_pff => xt_rsc_0_4_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_dp_inst : peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_4_i_qa_d => peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_dp_inst_xt_rsc_0_4_i_qa_d,
      xt_rsc_0_4_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_dp_inst_xt_rsc_0_4_i_qa_d_mxwt,
      xt_rsc_0_4_i_biwt => xt_rsc_0_4_i_biwt,
      xt_rsc_0_4_i_bdwt => xt_rsc_0_4_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_dp_inst_xt_rsc_0_4_i_qa_d <= xt_rsc_0_4_i_qa_d;
  xt_rsc_0_4_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_4_i_1_xt_rsc_0_4_wait_dp_inst_xt_rsc_0_4_i_qa_d_mxwt;

  xt_rsc_0_4_i_wea_d_pff <= xt_rsc_0_4_i_wea_d_core_sct_iff;
  xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_3_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_3_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_3_i_oswt : IN STD_LOGIC;
    xt_rsc_0_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_3_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_3_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_3_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_3_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_3_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_3_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_3_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_3_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_3_i_oswt : IN STD_LOGIC;
      xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_3_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_3_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_3_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_3_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_3_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_3_i_biwt : IN STD_LOGIC;
      xt_rsc_0_3_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_dp_inst_xt_rsc_0_3_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_dp_inst_xt_rsc_0_3_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_3_i_oswt => xt_rsc_0_3_i_oswt,
      xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_3_i_biwt => xt_rsc_0_3_i_biwt,
      xt_rsc_0_3_i_bdwt => xt_rsc_0_3_i_bdwt,
      xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_3_i_wea_d_core_sct_pff => xt_rsc_0_3_i_wea_d_core_sct_iff,
      xt_rsc_0_3_i_wea_d_core_psct_pff => xt_rsc_0_3_i_wea_d_core_psct_pff,
      xt_rsc_0_3_i_oswt_pff => xt_rsc_0_3_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_dp_inst : peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_3_i_qa_d => peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_dp_inst_xt_rsc_0_3_i_qa_d,
      xt_rsc_0_3_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_dp_inst_xt_rsc_0_3_i_qa_d_mxwt,
      xt_rsc_0_3_i_biwt => xt_rsc_0_3_i_biwt,
      xt_rsc_0_3_i_bdwt => xt_rsc_0_3_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_dp_inst_xt_rsc_0_3_i_qa_d <= xt_rsc_0_3_i_qa_d;
  xt_rsc_0_3_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_3_i_1_xt_rsc_0_3_wait_dp_inst_xt_rsc_0_3_i_qa_d_mxwt;

  xt_rsc_0_3_i_wea_d_pff <= xt_rsc_0_3_i_wea_d_core_sct_iff;
  xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_2_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_2_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_2_i_oswt : IN STD_LOGIC;
    xt_rsc_0_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_2_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_2_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_2_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_2_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_2_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_2_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_2_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_2_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_2_i_oswt : IN STD_LOGIC;
      xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_2_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_2_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_2_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_2_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_2_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_2_i_biwt : IN STD_LOGIC;
      xt_rsc_0_2_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_dp_inst_xt_rsc_0_2_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_dp_inst_xt_rsc_0_2_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_2_i_oswt => xt_rsc_0_2_i_oswt,
      xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_2_i_biwt => xt_rsc_0_2_i_biwt,
      xt_rsc_0_2_i_bdwt => xt_rsc_0_2_i_bdwt,
      xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_2_i_wea_d_core_sct_pff => xt_rsc_0_2_i_wea_d_core_sct_iff,
      xt_rsc_0_2_i_wea_d_core_psct_pff => xt_rsc_0_2_i_wea_d_core_psct_pff,
      xt_rsc_0_2_i_oswt_pff => xt_rsc_0_2_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_dp_inst : peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_2_i_qa_d => peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_dp_inst_xt_rsc_0_2_i_qa_d,
      xt_rsc_0_2_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_dp_inst_xt_rsc_0_2_i_qa_d_mxwt,
      xt_rsc_0_2_i_biwt => xt_rsc_0_2_i_biwt,
      xt_rsc_0_2_i_bdwt => xt_rsc_0_2_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_dp_inst_xt_rsc_0_2_i_qa_d <= xt_rsc_0_2_i_qa_d;
  xt_rsc_0_2_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_2_i_1_xt_rsc_0_2_wait_dp_inst_xt_rsc_0_2_i_qa_d_mxwt;

  xt_rsc_0_2_i_wea_d_pff <= xt_rsc_0_2_i_wea_d_core_sct_iff;
  xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_1_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_1_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_1_i_oswt : IN STD_LOGIC;
    xt_rsc_0_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_1_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_1_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_1_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_1_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_1_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_1_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_1_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_1_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_1_i_oswt : IN STD_LOGIC;
      xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_1_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_1_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_1_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_1_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_1_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_1_i_biwt : IN STD_LOGIC;
      xt_rsc_0_1_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_dp_inst_xt_rsc_0_1_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_dp_inst_xt_rsc_0_1_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_1_i_oswt => xt_rsc_0_1_i_oswt,
      xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_1_i_biwt => xt_rsc_0_1_i_biwt,
      xt_rsc_0_1_i_bdwt => xt_rsc_0_1_i_bdwt,
      xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_1_i_wea_d_core_sct_pff => xt_rsc_0_1_i_wea_d_core_sct_iff,
      xt_rsc_0_1_i_wea_d_core_psct_pff => xt_rsc_0_1_i_wea_d_core_psct_pff,
      xt_rsc_0_1_i_oswt_pff => xt_rsc_0_1_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_dp_inst : peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_1_i_qa_d => peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_dp_inst_xt_rsc_0_1_i_qa_d,
      xt_rsc_0_1_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_dp_inst_xt_rsc_0_1_i_qa_d_mxwt,
      xt_rsc_0_1_i_biwt => xt_rsc_0_1_i_biwt,
      xt_rsc_0_1_i_bdwt => xt_rsc_0_1_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_dp_inst_xt_rsc_0_1_i_qa_d <= xt_rsc_0_1_i_qa_d;
  xt_rsc_0_1_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_1_i_1_xt_rsc_0_1_wait_dp_inst_xt_rsc_0_1_i_qa_d_mxwt;

  xt_rsc_0_1_i_wea_d_pff <= xt_rsc_0_1_i_wea_d_core_sct_iff;
  xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core_xt_rsc_0_0_i_1
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core_xt_rsc_0_0_i_1 IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    core_wen : IN STD_LOGIC;
    xt_rsc_0_0_i_oswt : IN STD_LOGIC;
    core_wten : IN STD_LOGIC;
    xt_rsc_0_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
    xt_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_0_i_wea_d_core_psct_pff : IN STD_LOGIC;
    xt_rsc_0_0_i_oswt_pff : IN STD_LOGIC
  );
END peaseNTT_core_xt_rsc_0_0_i_1;

ARCHITECTURE v29 OF peaseNTT_core_xt_rsc_0_0_i_1 IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL xt_rsc_0_0_i_biwt : STD_LOGIC;
  SIGNAL xt_rsc_0_0_i_bdwt : STD_LOGIC;
  SIGNAL xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : STD_LOGIC;
  SIGNAL xt_rsc_0_0_i_wea_d_core_sct_iff : STD_LOGIC;

  COMPONENT peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_ctrl
    PORT(
      core_wen : IN STD_LOGIC;
      xt_rsc_0_0_i_oswt : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_0_i_biwt : OUT STD_LOGIC;
      xt_rsc_0_0_i_bdwt : OUT STD_LOGIC;
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct : OUT STD_LOGIC;
      xt_rsc_0_0_i_wea_d_core_sct_pff : OUT STD_LOGIC;
      xt_rsc_0_0_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_0_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_dp
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_0_i_biwt : IN STD_LOGIC;
      xt_rsc_0_0_i_bdwt : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_dp_inst_xt_rsc_0_0_i_qa_d :
      STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_dp_inst_xt_rsc_0_0_i_qa_d_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

BEGIN
  peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_ctrl_inst : peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_ctrl
    PORT MAP(
      core_wen => core_wen,
      xt_rsc_0_0_i_oswt => xt_rsc_0_0_i_oswt,
      core_wten => core_wten,
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct,
      xt_rsc_0_0_i_biwt => xt_rsc_0_0_i_biwt,
      xt_rsc_0_0_i_bdwt => xt_rsc_0_0_i_bdwt,
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct,
      xt_rsc_0_0_i_wea_d_core_sct_pff => xt_rsc_0_0_i_wea_d_core_sct_iff,
      xt_rsc_0_0_i_wea_d_core_psct_pff => xt_rsc_0_0_i_wea_d_core_psct_pff,
      xt_rsc_0_0_i_oswt_pff => xt_rsc_0_0_i_oswt_pff
    );
  peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_dp_inst : peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_dp
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_0_i_qa_d => peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_dp_inst_xt_rsc_0_0_i_qa_d,
      xt_rsc_0_0_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_dp_inst_xt_rsc_0_0_i_qa_d_mxwt,
      xt_rsc_0_0_i_biwt => xt_rsc_0_0_i_biwt,
      xt_rsc_0_0_i_bdwt => xt_rsc_0_0_i_bdwt
    );
  peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_dp_inst_xt_rsc_0_0_i_qa_d <= xt_rsc_0_0_i_qa_d;
  xt_rsc_0_0_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_0_i_1_xt_rsc_0_0_wait_dp_inst_xt_rsc_0_0_i_qa_d_mxwt;

  xt_rsc_0_0_i_wea_d_pff <= xt_rsc_0_0_i_wea_d_core_sct_iff;
  xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_sct;
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT_core
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT_core IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    xt_rsc_triosy_0_31_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_1_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_2_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_3_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_4_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_5_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_6_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_7_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_8_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_9_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_10_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_11_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_12_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_13_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_14_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_15_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_16_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_17_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_18_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_19_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_20_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_21_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_22_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_23_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_24_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_25_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_26_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_27_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_28_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_29_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_30_lz : OUT STD_LOGIC;
    xt_rsc_triosy_1_31_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_0_0_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_0_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_0_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_0_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_0_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_0_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_RID : OUT STD_LOGIC;
    twiddle_rsc_0_0_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_0_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_0_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_0_ARID : IN STD_LOGIC;
    twiddle_rsc_0_0_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_0_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_0_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_0_BID : OUT STD_LOGIC;
    twiddle_rsc_0_0_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_0_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_0_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_0_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_0_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_0_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_0_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_rsc_0_1_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_1_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_1_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_1_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_1_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_1_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_1_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_1_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_RID : OUT STD_LOGIC;
    twiddle_rsc_0_1_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_1_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_1_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_1_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_1_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_1_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_1_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_1_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_1_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_1_ARID : IN STD_LOGIC;
    twiddle_rsc_0_1_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_1_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_1_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_1_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_1_BID : OUT STD_LOGIC;
    twiddle_rsc_0_1_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_1_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_1_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_1_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_1_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_1_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_1_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_1_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_1_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_1_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_1_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_1_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_1_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_1_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_rsc_0_2_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_2_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_2_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_2_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_2_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_2_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_2_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_2_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_RID : OUT STD_LOGIC;
    twiddle_rsc_0_2_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_2_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_2_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_2_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_2_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_2_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_2_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_2_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_2_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_2_ARID : IN STD_LOGIC;
    twiddle_rsc_0_2_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_2_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_2_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_2_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_2_BID : OUT STD_LOGIC;
    twiddle_rsc_0_2_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_2_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_2_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_2_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_2_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_2_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_2_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_2_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_2_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_2_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_2_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_2_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_2_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_2_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_rsc_0_3_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_3_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_3_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_3_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_3_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_3_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_3_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_3_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_RID : OUT STD_LOGIC;
    twiddle_rsc_0_3_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_3_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_3_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_3_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_3_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_3_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_3_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_3_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_3_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_3_ARID : IN STD_LOGIC;
    twiddle_rsc_0_3_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_3_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_3_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_3_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_3_BID : OUT STD_LOGIC;
    twiddle_rsc_0_3_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_3_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_3_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_3_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_3_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_3_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_3_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_3_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_3_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_3_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_3_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_3_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_3_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_3_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_rsc_0_4_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_4_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_4_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_4_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_4_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_4_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_4_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_4_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_RID : OUT STD_LOGIC;
    twiddle_rsc_0_4_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_4_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_4_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_4_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_4_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_4_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_4_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_4_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_4_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_4_ARID : IN STD_LOGIC;
    twiddle_rsc_0_4_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_4_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_4_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_4_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_4_BID : OUT STD_LOGIC;
    twiddle_rsc_0_4_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_4_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_4_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_4_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_4_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_4_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_4_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_4_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_4_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_4_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_4_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_4_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_4_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_4_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_rsc_0_5_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_5_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_5_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_5_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_5_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_5_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_5_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_5_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_RID : OUT STD_LOGIC;
    twiddle_rsc_0_5_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_5_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_5_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_5_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_5_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_5_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_5_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_5_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_5_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_5_ARID : IN STD_LOGIC;
    twiddle_rsc_0_5_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_5_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_5_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_5_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_5_BID : OUT STD_LOGIC;
    twiddle_rsc_0_5_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_5_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_5_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_5_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_5_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_5_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_5_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_5_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_5_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_5_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_5_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_5_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_5_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_5_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_rsc_0_6_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_6_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_6_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_6_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_6_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_6_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_6_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_6_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_RID : OUT STD_LOGIC;
    twiddle_rsc_0_6_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_6_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_6_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_6_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_6_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_6_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_6_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_6_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_6_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_6_ARID : IN STD_LOGIC;
    twiddle_rsc_0_6_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_6_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_6_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_6_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_6_BID : OUT STD_LOGIC;
    twiddle_rsc_0_6_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_6_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_6_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_6_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_6_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_6_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_6_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_6_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_6_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_6_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_6_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_6_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_6_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_6_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_rsc_0_7_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_7_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_7_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_7_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_7_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_7_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_7_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_7_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_RID : OUT STD_LOGIC;
    twiddle_rsc_0_7_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_7_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_7_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_7_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_7_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_7_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_7_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_7_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_7_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_7_ARID : IN STD_LOGIC;
    twiddle_rsc_0_7_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_7_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_7_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_7_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_7_BID : OUT STD_LOGIC;
    twiddle_rsc_0_7_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_7_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_7_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_7_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_7_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_7_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_7_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_7_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_7_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_7_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_7_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_7_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_7_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_7_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_rsc_0_8_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_8_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_8_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_8_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_8_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_8_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_8_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_8_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_8_RID : OUT STD_LOGIC;
    twiddle_rsc_0_8_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_8_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_8_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_8_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_8_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_8_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_8_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_8_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_8_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_8_ARID : IN STD_LOGIC;
    twiddle_rsc_0_8_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_8_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_8_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_8_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_8_BID : OUT STD_LOGIC;
    twiddle_rsc_0_8_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_8_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_8_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_8_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_8_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_8_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_8_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_8_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_8_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_8_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_8_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_8_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_8_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_8_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_8_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_rsc_0_9_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_9_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_9_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_9_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_9_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_9_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_9_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_9_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_9_RID : OUT STD_LOGIC;
    twiddle_rsc_0_9_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_9_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_9_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_9_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_9_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_9_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_9_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_9_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_9_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_9_ARID : IN STD_LOGIC;
    twiddle_rsc_0_9_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_9_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_9_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_9_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_9_BID : OUT STD_LOGIC;
    twiddle_rsc_0_9_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_9_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_9_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_9_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_9_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_9_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_9_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_9_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_9_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_9_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_9_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_9_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_9_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_9_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_9_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_rsc_0_10_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_10_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_10_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_10_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_10_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_10_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_10_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_10_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_10_RID : OUT STD_LOGIC;
    twiddle_rsc_0_10_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_10_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_10_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_10_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_10_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_10_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_10_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_10_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_10_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_10_ARID : IN STD_LOGIC;
    twiddle_rsc_0_10_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_10_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_10_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_10_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_10_BID : OUT STD_LOGIC;
    twiddle_rsc_0_10_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_10_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_10_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_10_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_10_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_10_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_10_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_10_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_10_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_10_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_10_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_10_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_10_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_10_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_10_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_rsc_0_11_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_11_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_11_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_11_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_11_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_11_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_11_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_11_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_11_RID : OUT STD_LOGIC;
    twiddle_rsc_0_11_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_11_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_11_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_11_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_11_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_11_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_11_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_11_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_11_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_11_ARID : IN STD_LOGIC;
    twiddle_rsc_0_11_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_11_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_11_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_11_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_11_BID : OUT STD_LOGIC;
    twiddle_rsc_0_11_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_11_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_11_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_11_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_11_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_11_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_11_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_11_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_11_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_11_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_11_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_11_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_11_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_11_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_11_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_rsc_0_12_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_12_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_12_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_12_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_12_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_12_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_12_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_12_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_12_RID : OUT STD_LOGIC;
    twiddle_rsc_0_12_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_12_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_12_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_12_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_12_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_12_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_12_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_12_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_12_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_12_ARID : IN STD_LOGIC;
    twiddle_rsc_0_12_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_12_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_12_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_12_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_12_BID : OUT STD_LOGIC;
    twiddle_rsc_0_12_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_12_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_12_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_12_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_12_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_12_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_12_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_12_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_12_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_12_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_12_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_12_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_12_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_12_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_12_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_rsc_0_13_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_13_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_13_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_13_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_13_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_13_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_13_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_13_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_13_RID : OUT STD_LOGIC;
    twiddle_rsc_0_13_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_13_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_13_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_13_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_13_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_13_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_13_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_13_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_13_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_13_ARID : IN STD_LOGIC;
    twiddle_rsc_0_13_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_13_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_13_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_13_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_13_BID : OUT STD_LOGIC;
    twiddle_rsc_0_13_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_13_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_13_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_13_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_13_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_13_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_13_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_13_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_13_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_13_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_13_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_13_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_13_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_13_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_13_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_rsc_0_14_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_14_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_14_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_14_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_14_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_14_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_14_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_14_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_14_RID : OUT STD_LOGIC;
    twiddle_rsc_0_14_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_14_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_14_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_14_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_14_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_14_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_14_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_14_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_14_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_14_ARID : IN STD_LOGIC;
    twiddle_rsc_0_14_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_14_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_14_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_14_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_14_BID : OUT STD_LOGIC;
    twiddle_rsc_0_14_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_14_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_14_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_14_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_14_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_14_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_14_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_14_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_14_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_14_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_14_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_14_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_14_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_14_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_14_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_rsc_0_15_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_15_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_15_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_15_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_15_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_15_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_15_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_15_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_15_RID : OUT STD_LOGIC;
    twiddle_rsc_0_15_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_15_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_15_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_15_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_15_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_15_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_15_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_15_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_15_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_15_ARID : IN STD_LOGIC;
    twiddle_rsc_0_15_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_15_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_15_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_15_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_15_BID : OUT STD_LOGIC;
    twiddle_rsc_0_15_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_15_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_15_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_15_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_15_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_15_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_15_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_15_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_15_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_15_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_15_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_15_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_15_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_15_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_15_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_0_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_0_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_0_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_0_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_0_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_0_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_0_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_0_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_0_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_0_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_0_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_0_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_1_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_1_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_1_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_1_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_1_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_1_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_1_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_1_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_1_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_1_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_1_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_1_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_1_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_1_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_1_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_1_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_1_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_1_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_1_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_1_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_1_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_1_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_1_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_1_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_1_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_1_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_2_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_2_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_2_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_2_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_2_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_2_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_2_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_2_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_2_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_2_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_2_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_2_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_2_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_2_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_2_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_2_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_2_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_2_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_2_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_2_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_2_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_2_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_2_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_2_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_2_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_2_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_3_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_3_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_3_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_3_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_3_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_3_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_3_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_3_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_3_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_3_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_3_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_3_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_3_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_3_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_3_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_3_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_3_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_3_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_3_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_3_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_3_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_3_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_3_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_3_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_3_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_3_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_4_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_4_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_4_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_4_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_4_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_4_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_4_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_4_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_4_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_4_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_4_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_4_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_4_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_4_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_4_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_4_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_4_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_4_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_4_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_4_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_4_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_4_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_4_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_4_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_4_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_4_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_5_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_5_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_5_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_5_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_5_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_5_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_5_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_5_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_5_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_5_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_5_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_5_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_5_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_5_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_5_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_5_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_5_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_5_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_5_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_5_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_5_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_5_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_5_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_5_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_5_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_5_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_6_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_6_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_6_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_6_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_6_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_6_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_6_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_6_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_6_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_6_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_6_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_6_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_6_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_6_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_6_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_6_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_6_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_6_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_6_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_6_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_6_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_6_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_6_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_6_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_6_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_6_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_7_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_7_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_7_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_7_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_7_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_7_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_7_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_7_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_7_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_7_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_7_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_7_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_7_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_7_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_7_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_7_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_7_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_7_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_7_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_7_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_7_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_7_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_7_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_7_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_7_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_7_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_8_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_8_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_8_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_8_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_8_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_8_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_8_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_8_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_8_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_8_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_8_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_8_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_8_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_8_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_8_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_8_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_8_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_8_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_8_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_8_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_8_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_8_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_8_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_8_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_8_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_8_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_8_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_8_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_9_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_9_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_9_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_9_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_9_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_9_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_9_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_9_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_9_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_9_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_9_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_9_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_9_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_9_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_9_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_9_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_9_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_9_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_9_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_9_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_9_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_9_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_9_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_9_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_9_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_9_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_9_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_9_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_10_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_10_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_10_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_10_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_10_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_10_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_10_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_10_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_10_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_10_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_10_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_10_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_10_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_10_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_10_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_10_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_10_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_10_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_10_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_10_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_10_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_10_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_10_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_10_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_10_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_10_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_10_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_10_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_11_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_11_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_11_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_11_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_11_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_11_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_11_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_11_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_11_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_11_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_11_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_11_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_11_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_11_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_11_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_11_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_11_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_11_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_11_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_11_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_11_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_11_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_11_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_11_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_11_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_11_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_11_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_11_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_12_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_12_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_12_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_12_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_12_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_12_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_12_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_12_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_12_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_12_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_12_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_12_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_12_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_12_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_12_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_12_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_12_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_12_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_12_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_12_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_12_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_12_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_12_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_12_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_12_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_12_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_12_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_12_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_13_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_13_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_13_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_13_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_13_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_13_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_13_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_13_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_13_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_13_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_13_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_13_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_13_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_13_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_13_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_13_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_13_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_13_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_13_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_13_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_13_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_13_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_13_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_13_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_13_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_13_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_13_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_13_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_14_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_14_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_14_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_14_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_14_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_14_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_14_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_14_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_14_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_14_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_14_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_14_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_14_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_14_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_14_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_14_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_14_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_14_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_14_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_14_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_14_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_14_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_14_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_14_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_14_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_14_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_14_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_14_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_15_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_15_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_15_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_15_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_15_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_15_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_15_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_15_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_15_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_15_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_15_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_15_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_15_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_15_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_15_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_15_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_15_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_15_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_15_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_15_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_15_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_15_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_15_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_15_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_15_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_15_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_15_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_15_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    yt_rsc_0_0_i_clken_d : OUT STD_LOGIC;
    yt_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_16_i_clken_d : OUT STD_LOGIC;
    yt_rsc_0_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_0_i_clken_d : OUT STD_LOGIC;
    yt_rsc_1_0_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_1_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_2_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_3_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_4_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_5_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_6_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_7_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_8_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_9_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_10_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_11_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_12_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_13_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_14_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_15_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_16_i_clken_d : OUT STD_LOGIC;
    yt_rsc_1_16_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_17_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_18_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_19_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_20_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_21_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_22_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_23_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_24_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_25_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_26_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_27_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_28_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_29_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_30_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_31_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_1_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_0_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    xt_rsc_1_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
    yt_rsc_0_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
    yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    yt_rsc_0_1_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_2_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_3_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_4_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_5_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_6_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_7_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_8_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_9_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_10_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_11_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_12_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_13_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_14_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_15_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    yt_rsc_0_16_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_0_16_i_wea_d_pff : OUT STD_LOGIC;
    yt_rsc_1_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_1_0_i_wea_d_pff : OUT STD_LOGIC;
    yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
    yt_rsc_1_16_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    yt_rsc_1_16_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_1_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_1_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_2_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_2_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_3_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_3_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_4_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_4_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_5_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_5_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_6_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_6_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_7_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_7_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_8_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_8_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_9_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_9_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_10_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_10_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_11_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_11_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_12_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_12_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_13_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_13_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_14_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_14_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_15_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_15_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_16_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_16_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_17_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_18_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_19_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_20_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_21_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_22_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_23_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_24_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_25_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_26_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_27_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_28_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_29_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_30_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_0_31_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_0_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_1_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_1_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_2_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_2_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_3_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_3_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_4_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_4_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_5_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_5_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_6_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_6_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_7_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_7_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_8_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_8_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_9_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_9_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_10_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_10_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_11_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_11_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_12_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_12_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_13_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_13_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_14_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_14_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_15_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_15_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_16_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_17_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_18_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_19_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_20_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_21_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_22_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_23_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_24_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_25_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_26_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_27_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_28_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_29_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_30_i_wea_d_pff : OUT STD_LOGIC;
    xt_rsc_1_31_i_wea_d_pff : OUT STD_LOGIC
  );
END peaseNTT_core;

ARCHITECTURE v29 OF peaseNTT_core IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL core_wen : STD_LOGIC;
  SIGNAL p_rsci_idat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL core_wten : STD_LOGIC;
  SIGNAL xt_rsc_0_0_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_0_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_1_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_2_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_3_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_4_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_5_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_6_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_7_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_8_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_9_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_10_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_11_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_12_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_13_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_14_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_15_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_16_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_17_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_18_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_19_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_20_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_21_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_22_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_23_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_24_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_25_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_26_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_27_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_28_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_29_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_30_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_31_i_qa_d_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_0_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_1_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_1_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_2_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_2_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_3_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_3_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_4_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_4_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_5_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_5_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_6_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_6_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_7_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_7_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_8_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_8_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_9_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_9_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_10_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_10_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_11_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_11_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_12_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_12_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_13_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_13_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_14_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_14_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_rsc_0_15_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_rsc_0_15_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_0_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_1_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_1_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_2_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_2_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_3_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_3_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_4_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_4_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_5_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_5_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_6_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_6_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_7_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_7_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_8_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_8_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_9_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_9_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_10_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_10_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_11_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_11_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_12_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_12_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_13_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_13_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_14_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_14_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_15_i_wen_comp : STD_LOGIC;
  SIGNAL twiddle_h_rsc_0_15_i_s_din_mxwt : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_en : STD_LOGIC;
  SIGNAL mult_t_mul_cmp_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_1_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_2_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_3_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_4_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_5_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_6_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_7_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_8_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_9_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_10_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_11_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_12_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_13_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_14_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_15_z : STD_LOGIC_VECTOR (51 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_1_en : STD_LOGIC;
  SIGNAL mult_z_mul_cmp_1_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_2_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_3_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_4_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_5_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_6_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_7_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_8_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_9_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_10_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_11_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_12_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_13_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_14_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_15_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_16_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_17_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_18_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_19_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_20_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_21_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_22_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_23_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_24_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_25_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_26_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_27_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_28_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_29_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_30_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_31_z : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL twiddle_h_rsc_0_0_i_s_raddr_core_4 : STD_LOGIC;
  SIGNAL fsm_output : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL INNER_LOOP4_nor_tmp : STD_LOGIC;
  SIGNAL INNER_LOOP2_nor_tmp : STD_LOGIC;
  SIGNAL INNER_LOOP1_nor_tmp : STD_LOGIC;
  SIGNAL and_dcpl_144 : STD_LOGIC;
  SIGNAL and_dcpl_147 : STD_LOGIC;
  SIGNAL and_dcpl_149 : STD_LOGIC;
  SIGNAL and_dcpl_151 : STD_LOGIC;
  SIGNAL and_dcpl_153 : STD_LOGIC;
  SIGNAL and_dcpl_155 : STD_LOGIC;
  SIGNAL and_dcpl_157 : STD_LOGIC;
  SIGNAL and_dcpl_158 : STD_LOGIC;
  SIGNAL and_dcpl_159 : STD_LOGIC;
  SIGNAL and_dcpl_161 : STD_LOGIC;
  SIGNAL and_dcpl_163 : STD_LOGIC;
  SIGNAL and_dcpl_164 : STD_LOGIC;
  SIGNAL and_dcpl_165 : STD_LOGIC;
  SIGNAL and_dcpl_174 : STD_LOGIC;
  SIGNAL and_dcpl_175 : STD_LOGIC;
  SIGNAL and_dcpl_176 : STD_LOGIC;
  SIGNAL or_dcpl_29 : STD_LOGIC;
  SIGNAL or_tmp_804 : STD_LOGIC;
  SIGNAL or_tmp_806 : STD_LOGIC;
  SIGNAL or_tmp_812 : STD_LOGIC;
  SIGNAL or_tmp_814 : STD_LOGIC;
  SIGNAL or_tmp_827 : STD_LOGIC;
  SIGNAL or_tmp_835 : STD_LOGIC;
  SIGNAL or_tmp_888 : STD_LOGIC;
  SIGNAL or_tmp_895 : STD_LOGIC;
  SIGNAL and_252_cse : STD_LOGIC;
  SIGNAL and_253_cse : STD_LOGIC;
  SIGNAL and_655_cse : STD_LOGIC;
  SIGNAL and_656_cse : STD_LOGIC;
  SIGNAL and_1058_cse : STD_LOGIC;
  SIGNAL and_1059_cse : STD_LOGIC;
  SIGNAL and_1056_cse : STD_LOGIC;
  SIGNAL and_1057_cse : STD_LOGIC;
  SIGNAL and_1229_cse : STD_LOGIC;
  SIGNAL and_1230_cse : STD_LOGIC;
  SIGNAL and_1363_cse : STD_LOGIC;
  SIGNAL and_1364_cse : STD_LOGIC;
  SIGNAL and_1686_cse : STD_LOGIC;
  SIGNAL and_1695_cse : STD_LOGIC;
  SIGNAL and_1704_cse : STD_LOGIC;
  SIGNAL and_1929_cse : STD_LOGIC;
  SIGNAL and_1944_cse : STD_LOGIC;
  SIGNAL and_1948_cse : STD_LOGIC;
  SIGNAL and_1978_cse : STD_LOGIC;
  SIGNAL and_1994_cse : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_9_4_sva_2 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL INNER_LOOP4_r_9_4_sva_4_0 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL tmp_62_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_63_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_62_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_58_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_61_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_56_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_60_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_54_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_59_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_52_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_58_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_50_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_57_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_48_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_56_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_46_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_55_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_44_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_54_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_42_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_53_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_40_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_52_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_38_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_51_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_36_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_50_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_34_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_49_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_32_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_48_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP3_r_9_4_sva_4_0 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL tmp_126_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_47_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_46_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_45_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_44_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_43_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_42_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_41_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_40_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_39_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_38_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_37_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_36_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_35_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_100_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_34_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_98_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_33_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_96_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_32_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP2_r_9_4_sva_4_0 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL tmp_30_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_31_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_28_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_30_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_29_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_24_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_28_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_27_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_20_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_26_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_18_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_25_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_24_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_23_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_22_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_21_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_8_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_20_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_6_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_19_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_4_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_18_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_2_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_17_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_16_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_9_4_sva_2 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_9_4_sva_4_0 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL tmp_94_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_15_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_92_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_90_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_88_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_86_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_84_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_82_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_9_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_80_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_8_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_78_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_7_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_76_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_6_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_74_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_5_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_72_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_4_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_70_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_3_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_68_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_2_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_66_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_64_lpi_3_dfm_8 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_res_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly2_19_tw_asn_itm : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL c_1_sva : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_12 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_10 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_9 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_8 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_7 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_6 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_5 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_4 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_3 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_2 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_1 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_10 : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_9 : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_8 : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_7 : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_6 : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_5 : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_4 : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_3 : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_2 : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_1 : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm : STD_LOGIC;
  SIGNAL INNER_LOOP3_stage_0_12 : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_10 : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_9 : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_8 : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_7 : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_6 : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_5 : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_4 : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_3 : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_2 : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_1 : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_10 : STD_LOGIC;
  SIGNAL c_1_sva_1 : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_9 : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_8 : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_7 : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_6 : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_5 : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_4 : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_3 : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_2 : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_1 : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_191_itm_12 : STD_LOGIC;
  SIGNAL INNER_LOOP3_stage_0_13 : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_11 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_160_itm_12 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_13 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_11 : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4302_itm_1 : STD_LOGIC;
  SIGNAL INNER_LOOP2_stage_0_2 : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4377_itm_1 : STD_LOGIC;
  SIGNAL INNER_LOOP4_stage_0_2 : STD_LOGIC;
  SIGNAL INNER_LOOP3_stage_0 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0 : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_11 : STD_LOGIC;
  SIGNAL INNER_LOOP2_stage_0_12 : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_11 : STD_LOGIC;
  SIGNAL INNER_LOOP4_stage_0_12 : STD_LOGIC;
  SIGNAL operator_33_true_2_lshift_psp_2_0_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_33_true_3_lshift_psp_1_0_sva : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL INNER_LOOP4_stage_0 : STD_LOGIC;
  SIGNAL INNER_LOOP3_stage_0_2 : STD_LOGIC;
  SIGNAL INNER_LOOP3_stage_0_4 : STD_LOGIC;
  SIGNAL INNER_LOOP3_stage_0_3 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_3 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_2 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_4 : STD_LOGIC;
  SIGNAL INNER_LOOP2_stage_0_3 : STD_LOGIC;
  SIGNAL INNER_LOOP2_stage_0_4 : STD_LOGIC;
  SIGNAL INNER_LOOP4_stage_0_4 : STD_LOGIC;
  SIGNAL INNER_LOOP4_stage_0_3 : STD_LOGIC;
  SIGNAL INNER_LOOP3_stage_0_5 : STD_LOGIC;
  SIGNAL INNER_LOOP3_stage_0_6 : STD_LOGIC;
  SIGNAL INNER_LOOP3_stage_0_7 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_6 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_7 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_5 : STD_LOGIC;
  SIGNAL INNER_LOOP2_stage_0_6 : STD_LOGIC;
  SIGNAL INNER_LOOP2_stage_0_7 : STD_LOGIC;
  SIGNAL INNER_LOOP2_stage_0_5 : STD_LOGIC;
  SIGNAL INNER_LOOP4_stage_0_5 : STD_LOGIC;
  SIGNAL INNER_LOOP4_stage_0_6 : STD_LOGIC;
  SIGNAL INNER_LOOP4_stage_0_7 : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1 : STD_LOGIC;
  SIGNAL modulo_sub_base_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_1_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_2_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_3_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_4_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_5_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_6_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_7_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_8_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_9_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_10_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_11_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_12_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_13_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_14_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_15_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_15_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_14_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_13_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_12_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_11_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_10_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_9_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_8_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_7_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_6_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_5_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_4_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_3_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_2_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_1_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL modulo_sub_base_16_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_17_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_18_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_19_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_20_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_21_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_22_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_23_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_24_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_25_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_26_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_27_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_28_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_29_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_30_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_31_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP2_stage_0 : STD_LOGIC;
  SIGNAL mult_31_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_30_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_29_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_28_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_27_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_26_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_25_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_24_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_23_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_22_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_21_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_20_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_19_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_18_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_17_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_16_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL modulo_sub_base_32_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_33_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_34_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_35_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_36_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_37_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_38_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_39_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_40_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_41_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_42_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_43_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_44_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_45_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_46_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_47_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_47_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_46_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_45_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_44_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_43_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_42_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_41_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_40_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_39_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_38_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_37_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_36_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_35_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_34_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_33_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_32_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL modulo_sub_base_48_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_49_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_50_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_51_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_52_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_53_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_54_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_55_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_56_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_57_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_58_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_59_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_60_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_61_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_62_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_base_63_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_63_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_62_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_61_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_60_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_59_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_58_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_57_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_56_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_55_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_54_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_53_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_52_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_51_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_50_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_49_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL mult_48_slc_32_svs_st_1 : STD_LOGIC;
  SIGNAL modulo_add_base_63_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_62_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_61_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_60_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_59_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_58_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_57_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_56_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_55_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_54_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_53_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_52_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_51_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_50_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_49_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_48_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_63_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_62_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_61_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_60_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_59_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_58_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_57_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_56_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_55_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_54_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_53_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_52_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_51_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_50_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_49_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_48_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_47_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_46_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_45_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_44_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_43_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_42_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_41_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_40_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_39_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_38_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_37_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_36_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_35_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_34_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_33_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_32_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_47_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_46_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_45_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_44_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_43_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_42_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_41_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_40_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_39_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_38_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_37_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_36_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_35_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_34_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_33_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_32_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_31_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_30_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_29_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_28_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_27_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_26_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_25_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_24_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_23_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_22_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_21_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_20_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_19_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_18_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_17_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_16_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_31_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_30_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_29_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_28_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_27_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_26_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_25_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_15_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_14_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_13_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_12_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_11_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_10_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_9_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_8_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_7_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_6_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_5_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_4_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_3_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_2_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_1_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_base_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_15_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_9_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_8_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_7_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_6_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_5_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_4_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_3_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_2_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_res_sva_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_sva : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_15_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_15_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_15_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_14_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_14_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_14_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_13_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_13_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_13_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_12_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_12_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_12_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_11_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_11_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_11_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_10_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_10_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_10_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_9_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_9_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_9_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_8_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_8_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_8_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_7_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_7_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_7_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_6_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_6_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_6_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_5_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_5_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_5_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_4_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_4_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_4_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_3_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_3_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_3_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_2_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_2_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_2_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_1_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_1_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_1_and_ssc_3 : STD_LOGIC;
  SIGNAL butterFly1_and_ssc : STD_LOGIC;
  SIGNAL butterFly1_and_ssc_2 : STD_LOGIC;
  SIGNAL butterFly1_and_ssc_3 : STD_LOGIC;
  SIGNAL reg_yt_rsc_0_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_0_16_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_1_0_cgo_cse : STD_LOGIC;
  SIGNAL reg_yt_rsc_1_16_cgo_cse : STD_LOGIC;
  SIGNAL reg_xt_rsc_0_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_xt_rsc_0_16_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_xt_rsc_1_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_xt_rsc_1_16_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_0_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_1_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_2_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse : STD_LOGIC_VECTOR (4 DOWNTO
      0);
  SIGNAL reg_twiddle_rsc_0_3_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_4_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_5_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_6_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_7_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_8_i_oswt_cse : STD_LOGIC;
  SIGNAL reg_twiddle_rsc_0_0_i_s_raddr_core_3_0_cse : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL reg_xt_rsc_triosy_1_31_obj_iswt0_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_49_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_51_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_53_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_55_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_44_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_45_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_46_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_47_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_48_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_50_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_52_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_54_cse : STD_LOGIC;
  SIGNAL reg_ensig_cgo_17_cse : STD_LOGIC;
  SIGNAL reg_mult_15_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_14_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_13_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_12_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_11_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_10_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_9_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_8_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_7_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_6_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_5_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_4_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_3_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_2_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_1_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL reg_mult_z_asn_itm_1_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly2_7_tw_nor_cse : STD_LOGIC;
  SIGNAL butterFly2_7_tw_nor_1_cse : STD_LOGIC;
  SIGNAL butterFly2_7_tw_nor_2_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_or_9_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_or_10_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_or_11_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_or_12_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_41_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_42_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_43_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_37_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_38_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_39_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_30_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_31_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_32_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_or_3_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_40_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_36_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_and_29_cse : STD_LOGIC;
  SIGNAL c_or_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_or_1_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_tw_h_or_cse : STD_LOGIC;
  SIGNAL or_67_rmff : STD_LOGIC;
  SIGNAL or_166_rmff : STD_LOGIC;
  SIGNAL or_248_rmff : STD_LOGIC;
  SIGNAL butterFly1_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_1_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_1_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_2_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_2_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_3_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_3_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_4_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_4_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_5_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_5_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_6_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_6_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_7_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_7_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_8_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_8_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_9_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_9_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_10_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_10_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_11_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_11_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_12_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_12_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_13_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_13_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_14_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_14_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL butterFly1_15_and_4_rmff : STD_LOGIC;
  SIGNAL butterFly1_15_mux1h_2_rmff : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL or_347_rmff : STD_LOGIC;
  SIGNAL xt_rsc_0_0_i_wea_d_iff : STD_LOGIC;
  SIGNAL or_435_rmff : STD_LOGIC;
  SIGNAL or_429_rmff : STD_LOGIC;
  SIGNAL xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL or_436_rmff : STD_LOGIC;
  SIGNAL xt_rsc_0_1_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_2_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_3_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_4_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_5_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_6_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_7_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_8_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_9_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_10_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_11_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_12_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_13_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_14_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_15_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_16_i_wea_d_iff : STD_LOGIC;
  SIGNAL or_517_rmff : STD_LOGIC;
  SIGNAL or_512_rmff : STD_LOGIC;
  SIGNAL xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_17_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_18_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_19_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_20_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_21_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_22_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_23_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_24_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_25_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_26_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_27_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_28_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_29_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_30_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_0_31_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_0_i_wea_d_iff : STD_LOGIC;
  SIGNAL or_578_rmff : STD_LOGIC;
  SIGNAL xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL or_584_rmff : STD_LOGIC;
  SIGNAL xt_rsc_1_1_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_2_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_3_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_4_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_5_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_6_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_7_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_8_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_9_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_10_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_11_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_12_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_13_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_14_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_15_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_16_i_wea_d_iff : STD_LOGIC;
  SIGNAL or_660_rmff : STD_LOGIC;
  SIGNAL xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_17_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_18_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_19_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_20_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_21_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_22_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_23_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_24_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_25_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_26_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_27_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_28_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_29_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_30_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL xt_rsc_1_31_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg : STD_LOGIC;
  SIGNAL or_833_rmff : STD_LOGIC;
  SIGNAL or_956_rmff : STD_LOGIC;
  SIGNAL mult_4_t_mux1h_rmff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_65_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_1_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_a_mx0w2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_31_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_1_a_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_125_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_93_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_29_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_2_a_mx0w2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_3_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_91_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_27_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_121_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_5_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_89_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_25_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_4_a_mx0w2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_7_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_87_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_23_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_5_a_mx0w2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_12_a_mx0w3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_85_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_21_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_6_a_mx0w2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_11_a_mx0w3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_83_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_19_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_7_a_mx0w2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_10_a_mx0w3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_81_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_17_lpi_3_dfm_mx0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_8_a_mx0w2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_9_a_mx0w3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_9_a_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_9_a_mx0w2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_10_a_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_10_a_mx0w2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_11_a_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_11_a_mx0w2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_13_a_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_13_a_mx0w2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_14_a_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_14_a_mx0w2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_15_a_mx0w0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_15_a_mx0w2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_290_itm_11 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_321_itm_11 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL modulo_add_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_32_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_1_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_33_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_2_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_34_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_3_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_35_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_4_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_36_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_5_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_37_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_6_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_38_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_7_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_39_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_8_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_40_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_9_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_41_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_10_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_42_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_11_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_43_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_12_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_44_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_13_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_45_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_14_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_46_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_15_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_47_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_306_itm_11 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_337_itm_11 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_385_itm_10 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_416_itm_10 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_401_itm_10 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_432_itm_10 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_290_itm_11 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_321_itm_11 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL modulo_add_16_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_48_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_17_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_49_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_18_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_50_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_19_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_51_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_20_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_52_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_21_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_53_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_22_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_54_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_23_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_55_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_24_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_56_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_25_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_57_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_26_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_58_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_27_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_59_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_28_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_60_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_29_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_61_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_30_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_62_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_31_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_63_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_306_itm_11 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_337_itm_11 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL modulo_sub_16_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_48_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_17_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_49_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_18_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_50_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_19_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_51_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_20_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_52_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_21_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_53_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_22_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_54_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_23_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_55_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_24_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_56_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_25_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_57_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_26_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_58_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_27_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_59_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_28_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_60_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_29_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_61_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_30_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_62_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_31_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_63_qr_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_32 : STD_LOGIC_VECTOR (8 DOWNTO 0);
  SIGNAL z_out_33 : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL z_out_34 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_35 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_36 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_37 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_38 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_39 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_40 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_41 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_42 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_43 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_44 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_45 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_46 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_47 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_48 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_49 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_50 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_51 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_52 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_53 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_54 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_55 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_56 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_57 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_58 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_59 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_60 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_61 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_62 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_63 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_64 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_65 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_66 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_67 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_68 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_69 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_70 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_71 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_72 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_73 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_74 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_75 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_76 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_77 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_78 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_79 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_80 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_81 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_82 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_83 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_84 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_85 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_86 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_87 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_88 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_89 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_90 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_91 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_92 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_93 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_94 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_95 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_96 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_97 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_98 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_99 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_100 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_101 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_102 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_103 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_104 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_105 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_106 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_107 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_108 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL z_out_109 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL operator_20_false_acc_cse_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_33_true_return_8_4_sva : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL operator_33_true_1_lshift_psp_7_4_sva : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL INNER_LOOP1_stage_0_8 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_9 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_10 : STD_LOGIC;
  SIGNAL INNER_LOOP1_stage_0_11 : STD_LOGIC;
  SIGNAL tmp_64_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_64_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_64_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_64_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_64_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_64_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_64_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_66_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_66_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_66_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_66_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_66_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_66_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_66_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_68_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_68_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_68_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_68_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_68_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_68_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_68_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_2_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_70_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_70_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_70_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_70_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_70_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_70_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_70_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_3_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_72_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_72_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_72_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_72_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_72_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_72_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_72_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_4_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_74_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_74_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_74_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_74_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_74_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_74_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_74_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_5_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_76_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_76_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_76_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_76_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_76_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_76_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_76_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_6_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_78_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_78_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_78_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_78_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_78_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_78_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_78_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_7_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_80_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_80_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_80_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_80_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_80_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_80_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_80_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_8_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_82_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_82_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_82_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_82_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_82_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_82_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_82_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_9_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_84_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_84_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_84_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_84_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_84_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_84_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_84_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_86_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_86_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_86_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_86_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_86_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_86_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_86_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_88_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_88_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_88_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_88_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_88_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_88_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_88_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_90_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_90_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_90_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_90_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_90_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_90_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_90_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_92_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_92_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_92_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_92_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_92_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_92_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_92_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_94_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_94_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_94_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_94_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_94_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_94_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_94_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_15_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_1_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_2_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_2_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_2_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_2_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_3_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_3_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_3_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_3_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_4_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_4_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_4_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_4_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_5_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_5_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_5_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_5_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_6_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_6_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_6_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_6_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_7_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_7_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_7_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_7_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_8_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_8_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_8_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_8_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_9_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_9_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_9_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_9_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_10_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_11_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_12_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_13_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_14_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_15_z_asn_itm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_15_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_15_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_15_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_1 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_2 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_3 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_4 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_5 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_6 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_7 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_8 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_9 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_1 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_2 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_3 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_4 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_5 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_6 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_7 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_8 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_9 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP2_stage_0_8 : STD_LOGIC;
  SIGNAL INNER_LOOP2_stage_0_9 : STD_LOGIC;
  SIGNAL INNER_LOOP2_stage_0_10 : STD_LOGIC;
  SIGNAL INNER_LOOP2_stage_0_11 : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4302_itm : STD_LOGIC;
  SIGNAL tmp_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_16_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_2_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_2_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_2_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_2_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_2_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_2_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_2_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_17_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_4_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_4_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_4_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_4_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_4_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_4_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_4_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_18_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_6_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_6_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_6_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_6_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_6_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_6_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_6_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_19_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_8_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_8_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_8_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_8_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_8_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_8_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_8_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_20_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_10_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_21_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_12_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_22_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_14_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_23_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_16_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_24_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_18_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_18_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_18_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_18_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_18_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_18_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_18_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_25_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_20_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_20_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_20_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_20_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_20_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_20_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_20_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_26_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_22_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_27_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_24_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_24_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_24_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_24_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_24_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_24_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_24_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_28_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_26_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_29_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_28_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_28_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_28_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_28_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_28_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_28_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_28_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_30_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_30_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_30_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_30_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_30_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_30_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_30_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_30_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_31_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_16_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_16_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_16_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_17_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_17_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_17_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_18_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_18_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_18_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_19_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_19_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_19_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_20_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_20_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_20_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_21_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_21_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_21_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_22_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_22_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_22_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_23_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_23_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_23_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_24_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_24_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_24_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_25_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_25_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_25_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_26_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_26_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_26_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_27_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_27_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_27_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_28_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_28_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_28_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_29_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_29_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_29_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_30_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_30_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_30_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_31_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_31_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_31_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_1 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_2 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_3 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_4 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_5 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_6 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_7 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_8 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_9 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_10 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_1 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_2 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_3 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_4 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_5 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_6 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_7 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_8 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_9 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_10 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP3_stage_0_8 : STD_LOGIC;
  SIGNAL INNER_LOOP3_stage_0_9 : STD_LOGIC;
  SIGNAL INNER_LOOP3_stage_0_10 : STD_LOGIC;
  SIGNAL INNER_LOOP3_stage_0_11 : STD_LOGIC;
  SIGNAL tmp_96_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_96_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_96_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_96_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_96_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_96_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_96_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_32_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_98_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_98_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_98_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_98_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_98_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_98_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_98_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_33_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_100_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_100_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_100_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_100_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_100_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_100_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_100_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_34_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_102_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_35_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_104_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_36_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_106_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_37_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_108_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_38_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_110_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_39_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_112_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_40_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_114_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_41_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_116_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_42_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_118_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_43_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_120_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_44_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_122_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_45_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_124_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_46_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_lpi_3_dfm_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_126_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly2_15_tw_equal_tmp_1 : STD_LOGIC;
  SIGNAL butterFly2_15_tw_equal_tmp_3_1 : STD_LOGIC;
  SIGNAL butterFly2_15_tw_equal_tmp_5_1 : STD_LOGIC;
  SIGNAL butterFly2_15_tw_equal_tmp_6_1 : STD_LOGIC;
  SIGNAL butterFly2_15_tw_equal_tmp_7_1 : STD_LOGIC;
  SIGNAL mult_47_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_32_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_32_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_32_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_33_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_33_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_33_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_34_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_34_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_34_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_35_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_35_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_35_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_36_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_36_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_36_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_37_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_37_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_37_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_38_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_38_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_38_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_39_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_39_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_39_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_40_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_40_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_40_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_41_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_41_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_41_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_42_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_42_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_42_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_43_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_43_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_43_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_44_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_44_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_44_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_45_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_45_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_45_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_46_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_46_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_46_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_47_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_47_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_47_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_1 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_2 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_3 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_4 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_5 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_6 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_7 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_8 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_9 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_1 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_2 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_3 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_4 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_5 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_6 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_7 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_8 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_9 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP4_stage_0_8 : STD_LOGIC;
  SIGNAL INNER_LOOP4_stage_0_9 : STD_LOGIC;
  SIGNAL INNER_LOOP4_stage_0_10 : STD_LOGIC;
  SIGNAL INNER_LOOP4_stage_0_11 : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4377_itm : STD_LOGIC;
  SIGNAL tmp_32_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_32_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_32_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_32_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_32_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_32_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_48_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_34_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_34_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_34_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_34_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_34_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_34_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_49_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_36_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_36_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_36_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_36_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_36_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_36_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_50_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_38_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_38_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_38_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_38_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_38_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_38_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_51_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_40_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_40_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_40_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_40_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_40_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_40_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_52_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_42_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_42_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_42_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_42_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_42_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_42_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_53_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_44_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_44_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_44_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_44_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_44_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_44_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_54_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_46_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_46_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_46_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_46_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_46_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_46_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_55_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_48_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_48_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_48_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_48_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_48_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_48_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_56_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_50_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_50_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_50_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_50_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_50_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_50_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_57_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_52_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_52_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_52_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_52_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_52_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_52_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_58_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_54_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_54_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_54_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_54_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_54_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_54_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_59_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_56_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_56_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_56_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_56_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_56_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_56_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_60_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_58_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_58_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_58_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_58_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_58_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_58_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_61_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_60_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_62_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_lpi_3_dfm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_lpi_3_dfm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_lpi_3_dfm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_lpi_3_dfm_5 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_lpi_3_dfm_6 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL tmp_62_lpi_3_dfm_7 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_63_res_sva_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_48_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_48_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_48_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_49_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_49_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_49_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_50_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_50_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_50_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_51_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_51_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_51_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_52_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_52_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_52_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_53_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_53_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_53_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_54_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_54_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_54_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_55_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_55_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_55_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_56_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_56_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_56_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_57_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_57_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_57_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_58_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_58_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_58_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_59_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_59_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_59_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_60_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_60_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_60_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_61_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_61_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_61_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_62_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_62_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_62_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_63_z_asn_itm_2 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_63_z_asn_itm_3 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_63_z_asn_itm_4 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_1 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_2 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_3 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_4 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_5 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_6 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_7 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_8 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_9 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_10 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_1 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_2 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_3 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_4 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_5 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_6 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_7 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_8 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_9 : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_10 : STD_LOGIC_VECTOR (3
      DOWNTO 0);
  SIGNAL operator_33_true_3_lshift_psp_1_0_sva_mx0w2 : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL operator_20_false_acc_cse_sva_mx0w0 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL INNER_LOOP1_tw_and_psp_sva_1 : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL modulo_add_qelse_and_cse : STD_LOGIC;
  SIGNAL butterFly1_and_cse : STD_LOGIC;
  SIGNAL mult_15_if_and_cse : STD_LOGIC;
  SIGNAL and_1665_cse : STD_LOGIC;
  SIGNAL mult_15_z_and_cse : STD_LOGIC;
  SIGNAL mult_15_z_and_cse_1 : STD_LOGIC;
  SIGNAL mult_15_z_and_1_cse : STD_LOGIC;
  SIGNAL mult_15_z_and_2_cse : STD_LOGIC;
  SIGNAL mult_15_z_and_3_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_and_20_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_and_23_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_and_26_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_and_29_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_and_7_cse : STD_LOGIC;
  SIGNAL modulo_add_16_qelse_and_cse : STD_LOGIC;
  SIGNAL butterFly1_31_and_cse : STD_LOGIC;
  SIGNAL mult_31_if_and_cse : STD_LOGIC;
  SIGNAL and_1666_cse : STD_LOGIC;
  SIGNAL mult_31_z_and_cse : STD_LOGIC;
  SIGNAL mult_31_z_and_1_cse : STD_LOGIC;
  SIGNAL mult_31_z_and_2_cse : STD_LOGIC;
  SIGNAL butterFly1_31_f1_and_4_cse : STD_LOGIC;
  SIGNAL butterFly1_31_f1_and_5_cse : STD_LOGIC;
  SIGNAL butterFly1_31_f1_and_6_cse : STD_LOGIC;
  SIGNAL butterFly1_31_f1_and_7_cse : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_and_3_cse : STD_LOGIC;
  SIGNAL INNER_LOOP2_r_and_4_cse : STD_LOGIC;
  SIGNAL modulo_add_32_qelse_and_cse : STD_LOGIC;
  SIGNAL butterFly2_and_cse : STD_LOGIC;
  SIGNAL mult_47_if_and_cse : STD_LOGIC;
  SIGNAL butterFly2_15_tw_and_cse : STD_LOGIC;
  SIGNAL mult_47_z_and_cse : STD_LOGIC;
  SIGNAL mult_47_z_and_1_cse : STD_LOGIC;
  SIGNAL mult_47_z_and_2_cse : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_and_19_cse : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_and_22_cse : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_and_25_cse : STD_LOGIC;
  SIGNAL INNER_LOOP3_r_and_28_cse : STD_LOGIC;
  SIGNAL modulo_add_48_qelse_and_cse : STD_LOGIC;
  SIGNAL butterFly2_31_and_cse : STD_LOGIC;
  SIGNAL mult_63_if_and_cse : STD_LOGIC;
  SIGNAL mult_63_z_and_cse : STD_LOGIC;
  SIGNAL mult_63_z_and_1_cse : STD_LOGIC;
  SIGNAL mult_63_z_and_2_cse : STD_LOGIC;
  SIGNAL butterFly2_31_f1_and_4_cse : STD_LOGIC;
  SIGNAL butterFly2_31_f1_and_5_cse : STD_LOGIC;
  SIGNAL butterFly2_31_f1_and_6_cse : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_and_3_cse : STD_LOGIC;
  SIGNAL INNER_LOOP4_r_and_4_cse : STD_LOGIC;
  SIGNAL INNER_LOOP1_r_INNER_LOOP1_r_and_2_cse : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL INNER_LOOP1_r_INNER_LOOP1_r_and_6_cse : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL INNER_LOOP4_INNER_LOOP4_and_1_cse : STD_LOGIC;
  SIGNAL INNER_LOOP3_INNER_LOOP3_and_1_cse : STD_LOGIC;
  SIGNAL z_out_32_1 : STD_LOGIC;
  SIGNAL z_out_1_32 : STD_LOGIC;
  SIGNAL z_out_2_32 : STD_LOGIC;
  SIGNAL z_out_3_32 : STD_LOGIC;
  SIGNAL z_out_4_32 : STD_LOGIC;
  SIGNAL z_out_5_32 : STD_LOGIC;
  SIGNAL z_out_6_32 : STD_LOGIC;
  SIGNAL z_out_7_32 : STD_LOGIC;
  SIGNAL z_out_8_32 : STD_LOGIC;
  SIGNAL z_out_9_32 : STD_LOGIC;
  SIGNAL z_out_10_32 : STD_LOGIC;
  SIGNAL z_out_11_32 : STD_LOGIC;
  SIGNAL z_out_12_32 : STD_LOGIC;
  SIGNAL z_out_13_32 : STD_LOGIC;
  SIGNAL z_out_14_32 : STD_LOGIC;
  SIGNAL z_out_15_32 : STD_LOGIC;
  SIGNAL z_out_16_32 : STD_LOGIC;
  SIGNAL z_out_17_32 : STD_LOGIC;
  SIGNAL z_out_18_32 : STD_LOGIC;
  SIGNAL z_out_19_32 : STD_LOGIC;
  SIGNAL z_out_20_32 : STD_LOGIC;
  SIGNAL z_out_21_32 : STD_LOGIC;
  SIGNAL z_out_22_32 : STD_LOGIC;
  SIGNAL z_out_23_32 : STD_LOGIC;
  SIGNAL z_out_24_32 : STD_LOGIC;
  SIGNAL z_out_25_32 : STD_LOGIC;
  SIGNAL z_out_26_32 : STD_LOGIC;
  SIGNAL z_out_27_32 : STD_LOGIC;
  SIGNAL z_out_28_32 : STD_LOGIC;
  SIGNAL z_out_29_32 : STD_LOGIC;
  SIGNAL z_out_30_32 : STD_LOGIC;
  SIGNAL z_out_31_32 : STD_LOGIC;
  SIGNAL butterFly1_10_mux_7_cse : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL INNER_LOOP2_tw_and_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL mult_4_t_and_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_1_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_2_nl : STD_LOGIC;
  SIGNAL mult_4_t_and_3_nl : STD_LOGIC;
  SIGNAL nor_4_nl : STD_LOGIC;
  SIGNAL modulo_add_20_qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_21_qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_22_qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_23_qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_24_qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_25_qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_26_qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_27_qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_28_qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_29_qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_30_qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_31_qif_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_31_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_30_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_29_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_28_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_27_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_26_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_25_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_24_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_23_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_22_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_21_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_20_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_19_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_18_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_17_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_16_if_acc_1_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly2_21_tw_butterFly2_21_tw_or_nl : STD_LOGIC;
  SIGNAL mult_22_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_21_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_20_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_19_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_18_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_17_if_acc_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_1_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_1_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_2_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_2_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_3_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_3_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_4_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_4_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_5_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_5_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_6_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_6_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_7_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_7_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_8_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_8_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_9_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_9_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_10_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_10_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_11_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_11_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_12_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_12_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_13_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_13_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_14_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_14_and_1_nl : STD_LOGIC;
  SIGNAL butterFly1_15_mux_nl : STD_LOGIC;
  SIGNAL butterFly1_15_and_1_nl : STD_LOGIC;
  SIGNAL acc_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_1_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_1_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_2_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_2_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_3_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_3_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_4_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_4_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_5_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_5_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_6_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_6_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_7_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_7_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_8_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_8_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_9_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_9_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_10_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_10_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_11_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_11_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_12_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_12_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_13_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_13_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_14_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_14_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_15_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL modulo_add_15_mux1h_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_16_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_15_if_mux1h_4_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_17_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_14_if_mux1h_4_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_18_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_13_if_mux1h_4_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_19_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_12_if_mux1h_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_20_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_11_if_mux1h_4_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_21_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_10_if_mux1h_4_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_22_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_9_if_mux1h_4_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_23_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_8_if_mux1h_4_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_24_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_7_if_mux1h_4_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_25_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_6_if_mux1h_4_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_26_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_5_if_mux1h_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_27_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_4_if_mux1h_4_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_28_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_3_if_mux1h_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_29_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_2_if_mux1h_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_30_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_1_if_mux1h_4_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_31_nl : STD_LOGIC_VECTOR (33 DOWNTO 0);
  SIGNAL mult_if_mux1h_6_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL operator_20_false_1_mux_2_nl : STD_LOGIC_VECTOR (4 DOWNTO 0);
  SIGNAL acc_33_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_40_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_34_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_41_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_35_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_42_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_63_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_37_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_63_qif_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_62_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_39_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_62_qif_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_62_qif_mux_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_61_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_41_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_61_qif_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_61_qif_mux_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_60_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_43_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_60_qif_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_60_qif_mux_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_59_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_45_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_59_qif_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_59_qif_mux_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_58_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_47_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_58_qif_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_58_qif_mux_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_57_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_16_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_50_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_12_if_mux1h_7_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_17_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_52_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_47_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_18_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_54_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_54_qif_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_54_qif_mux_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_19_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_56_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_46_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_20_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_58_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_45_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_21_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_60_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_44_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_22_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_62_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_43_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_sub_23_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_56_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_24_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_55_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_25_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_54_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_26_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_53_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_27_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_52_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_28_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_51_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_29_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_50_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_30_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_48_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_31_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL modulo_sub_49_qif_mux_2_nl : STD_LOGIC_VECTOR (30 DOWNTO 0);
  SIGNAL acc_81_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_57_qif_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_57_qif_mux_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_82_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_55_qif_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_55_qif_mux_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_83_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_56_qif_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL modulo_add_56_qif_mux_3_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL butterFly1_10_mux_8_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_85_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL butterFly1_10_mux_10_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_86_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_87_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_1_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_88_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_2_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_89_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_3_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_90_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_4_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_91_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_5_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_92_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_6_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_93_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_7_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_94_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_8_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_95_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_9_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_96_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_10_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_97_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_11_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_98_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_12_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_99_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_13_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_100_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_14_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_101_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_15_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_102_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_5_if_mux1h_7_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_103_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_3_if_mux1h_7_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_104_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_if_mux1h_7_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_105_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_16_if_mux_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_106_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL mult_2_if_mux1h_7_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_107_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_51_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL acc_108_nl : STD_LOGIC_VECTOR (32 DOWNTO 0);
  SIGNAL modulo_add_53_qif_mux1h_2_nl : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_rsci_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL p_rsci_idat_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_1_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_1_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_1_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_2_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_2_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_2_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_3_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_3_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_3_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_4_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_4_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_4_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_5_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_5_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_5_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_6_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_6_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_6_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_7_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_7_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_7_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_8_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_8_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_8_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_9_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_9_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_9_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_10_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_10_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_10_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_11_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_11_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_11_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_12_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_12_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_12_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_13_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_13_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_13_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_14_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_14_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_14_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_t_mul_cmp_15_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_15_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_t_mul_cmp_15_z_1 : STD_LOGIC_VECTOR (51 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_1_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_1_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_1_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_2_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_2_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_2_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_3_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_3_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_3_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_4_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_4_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_4_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_5_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_5_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_5_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_6_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_6_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_6_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_7_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_7_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_7_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_8_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_8_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_8_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_9_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_9_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_9_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_10_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_10_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_10_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_11_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_11_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_11_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_12_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_12_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_12_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_13_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_13_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_13_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_14_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_14_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_14_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_15_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_15_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_15_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_16_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_16_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_16_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_17_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_17_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_17_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_18_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_18_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_18_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_19_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_19_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_19_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_20_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_20_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_20_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_21_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_21_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_21_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_22_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_22_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_22_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_23_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_23_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_23_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_24_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_24_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_24_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_25_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_25_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_25_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_26_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_26_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_26_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_27_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_27_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_27_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_28_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_28_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_28_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_29_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_29_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_29_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_30_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_30_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_30_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL mult_z_mul_cmp_31_a : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_31_b : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL mult_z_mul_cmp_31_z_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL operator_33_true_3_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL operator_33_true_3_lshift_rg_s : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL operator_33_true_3_lshift_rg_z : STD_LOGIC_VECTOR (1 DOWNTO 0);

  SIGNAL operator_33_true_1_lshift_rg_a : STD_LOGIC_VECTOR (0 DOWNTO 0);
  SIGNAL operator_33_true_1_lshift_rg_s : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL operator_33_true_1_lshift_rg_z : STD_LOGIC_VECTOR (8 DOWNTO 0);

  COMPONENT peaseNTT_core_wait_dp
    PORT(
      yt_rsc_0_0_cgo_iro : IN STD_LOGIC;
      yt_rsc_0_0_i_clken_d : OUT STD_LOGIC;
      yt_rsc_0_16_cgo_iro : IN STD_LOGIC;
      yt_rsc_0_16_i_clken_d : OUT STD_LOGIC;
      yt_rsc_1_0_cgo_iro : IN STD_LOGIC;
      yt_rsc_1_0_i_clken_d : OUT STD_LOGIC;
      yt_rsc_1_16_cgo_iro : IN STD_LOGIC;
      yt_rsc_1_16_i_clken_d : OUT STD_LOGIC;
      ensig_cgo_iro : IN STD_LOGIC;
      ensig_cgo_iro_17 : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      yt_rsc_0_0_cgo : IN STD_LOGIC;
      yt_rsc_0_16_cgo : IN STD_LOGIC;
      yt_rsc_1_0_cgo : IN STD_LOGIC;
      yt_rsc_1_16_cgo : IN STD_LOGIC;
      ensig_cgo : IN STD_LOGIC;
      mult_t_mul_cmp_en : OUT STD_LOGIC;
      ensig_cgo_17 : IN STD_LOGIC;
      mult_z_mul_cmp_1_en : OUT STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_0_0_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      xt_rsc_0_0_i_oswt : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_0_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_0_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_0_i_1_inst_xt_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_0_i_1_inst_xt_rsc_0_0_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_1_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_1_i_oswt : IN STD_LOGIC;
      xt_rsc_0_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_1_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_1_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_1_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_1_i_1_inst_xt_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_1_i_1_inst_xt_rsc_0_1_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_2_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_2_i_oswt : IN STD_LOGIC;
      xt_rsc_0_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_2_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_2_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_2_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_2_i_1_inst_xt_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_2_i_1_inst_xt_rsc_0_2_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_3_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_3_i_oswt : IN STD_LOGIC;
      xt_rsc_0_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_3_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_3_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_3_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_3_i_1_inst_xt_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_3_i_1_inst_xt_rsc_0_3_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_4_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_4_i_oswt : IN STD_LOGIC;
      xt_rsc_0_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_4_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_4_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_4_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_4_i_1_inst_xt_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_4_i_1_inst_xt_rsc_0_4_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_5_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_5_i_oswt : IN STD_LOGIC;
      xt_rsc_0_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_5_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_5_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_5_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_5_i_1_inst_xt_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_5_i_1_inst_xt_rsc_0_5_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_6_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_6_i_oswt : IN STD_LOGIC;
      xt_rsc_0_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_6_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_6_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_6_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_6_i_1_inst_xt_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_6_i_1_inst_xt_rsc_0_6_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_7_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_7_i_oswt : IN STD_LOGIC;
      xt_rsc_0_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_7_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_7_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_7_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_7_i_1_inst_xt_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_7_i_1_inst_xt_rsc_0_7_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_8_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_8_i_oswt : IN STD_LOGIC;
      xt_rsc_0_8_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_8_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_8_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_8_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_8_i_1_inst_xt_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_8_i_1_inst_xt_rsc_0_8_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_9_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_9_i_oswt : IN STD_LOGIC;
      xt_rsc_0_9_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_9_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_9_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_9_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_9_i_1_inst_xt_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_9_i_1_inst_xt_rsc_0_9_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_10_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_10_i_oswt : IN STD_LOGIC;
      xt_rsc_0_10_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_10_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_10_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_10_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_10_i_1_inst_xt_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_10_i_1_inst_xt_rsc_0_10_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_11_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_11_i_oswt : IN STD_LOGIC;
      xt_rsc_0_11_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_11_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_11_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_11_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_11_i_1_inst_xt_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_11_i_1_inst_xt_rsc_0_11_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_12_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_12_i_oswt : IN STD_LOGIC;
      xt_rsc_0_12_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_12_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_12_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_12_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_12_i_1_inst_xt_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_12_i_1_inst_xt_rsc_0_12_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_13_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_13_i_oswt : IN STD_LOGIC;
      xt_rsc_0_13_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_13_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_13_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_13_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_13_i_1_inst_xt_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_13_i_1_inst_xt_rsc_0_13_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_14_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_14_i_oswt : IN STD_LOGIC;
      xt_rsc_0_14_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_14_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_14_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_14_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_14_i_1_inst_xt_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_14_i_1_inst_xt_rsc_0_14_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_15_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_15_i_oswt : IN STD_LOGIC;
      xt_rsc_0_15_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_15_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_15_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_15_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_15_i_1_inst_xt_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_15_i_1_inst_xt_rsc_0_15_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_16_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_16_i_oswt : IN STD_LOGIC;
      xt_rsc_0_16_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_16_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_16_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_16_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_16_i_1_inst_xt_rsc_0_16_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_16_i_1_inst_xt_rsc_0_16_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_17_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_17_i_oswt : IN STD_LOGIC;
      xt_rsc_0_17_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_17_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_17_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_17_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_17_i_1_inst_xt_rsc_0_17_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_17_i_1_inst_xt_rsc_0_17_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_18_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_18_i_oswt : IN STD_LOGIC;
      xt_rsc_0_18_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_18_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_18_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_18_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_18_i_1_inst_xt_rsc_0_18_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_18_i_1_inst_xt_rsc_0_18_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_19_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_19_i_oswt : IN STD_LOGIC;
      xt_rsc_0_19_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_19_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_19_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_19_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_19_i_1_inst_xt_rsc_0_19_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_19_i_1_inst_xt_rsc_0_19_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_20_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_20_i_oswt : IN STD_LOGIC;
      xt_rsc_0_20_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_20_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_20_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_20_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_20_i_1_inst_xt_rsc_0_20_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_20_i_1_inst_xt_rsc_0_20_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_21_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_21_i_oswt : IN STD_LOGIC;
      xt_rsc_0_21_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_21_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_21_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_21_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_21_i_1_inst_xt_rsc_0_21_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_21_i_1_inst_xt_rsc_0_21_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_22_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_22_i_oswt : IN STD_LOGIC;
      xt_rsc_0_22_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_22_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_22_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_22_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_22_i_1_inst_xt_rsc_0_22_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_22_i_1_inst_xt_rsc_0_22_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_23_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_23_i_oswt : IN STD_LOGIC;
      xt_rsc_0_23_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_23_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_23_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_23_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_23_i_1_inst_xt_rsc_0_23_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_23_i_1_inst_xt_rsc_0_23_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_24_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_24_i_oswt : IN STD_LOGIC;
      xt_rsc_0_24_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_24_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_24_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_24_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_24_i_1_inst_xt_rsc_0_24_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_24_i_1_inst_xt_rsc_0_24_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_25_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_25_i_oswt : IN STD_LOGIC;
      xt_rsc_0_25_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_25_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_25_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_25_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_25_i_1_inst_xt_rsc_0_25_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_25_i_1_inst_xt_rsc_0_25_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_26_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_26_i_oswt : IN STD_LOGIC;
      xt_rsc_0_26_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_26_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_26_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_26_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_26_i_1_inst_xt_rsc_0_26_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_26_i_1_inst_xt_rsc_0_26_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_27_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_27_i_oswt : IN STD_LOGIC;
      xt_rsc_0_27_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_27_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_27_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_27_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_27_i_1_inst_xt_rsc_0_27_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_27_i_1_inst_xt_rsc_0_27_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_28_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_28_i_oswt : IN STD_LOGIC;
      xt_rsc_0_28_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_28_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_28_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_28_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_28_i_1_inst_xt_rsc_0_28_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_28_i_1_inst_xt_rsc_0_28_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_29_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_29_i_oswt : IN STD_LOGIC;
      xt_rsc_0_29_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_29_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_29_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_29_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_29_i_1_inst_xt_rsc_0_29_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_29_i_1_inst_xt_rsc_0_29_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_30_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_30_i_oswt : IN STD_LOGIC;
      xt_rsc_0_30_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_30_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_30_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_30_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_30_i_1_inst_xt_rsc_0_30_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_30_i_1_inst_xt_rsc_0_30_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_0_31_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_0_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_0_31_i_oswt : IN STD_LOGIC;
      xt_rsc_0_31_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_0_31_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_31_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_0_31_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_0_31_i_1_inst_xt_rsc_0_31_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_0_31_i_1_inst_xt_rsc_0_31_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_0_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_0_i_oswt : IN STD_LOGIC;
      xt_rsc_1_0_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_0_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_0_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_0_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_0_i_1_inst_xt_rsc_1_0_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_0_i_1_inst_xt_rsc_1_0_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_1_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_1_i_oswt : IN STD_LOGIC;
      xt_rsc_1_1_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_1_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_1_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_1_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_1_i_1_inst_xt_rsc_1_1_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_1_i_1_inst_xt_rsc_1_1_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_2_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_2_i_oswt : IN STD_LOGIC;
      xt_rsc_1_2_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_2_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_2_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_2_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_2_i_1_inst_xt_rsc_1_2_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_2_i_1_inst_xt_rsc_1_2_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_3_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_3_i_oswt : IN STD_LOGIC;
      xt_rsc_1_3_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_3_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_3_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_3_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_3_i_1_inst_xt_rsc_1_3_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_3_i_1_inst_xt_rsc_1_3_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_4_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_4_i_oswt : IN STD_LOGIC;
      xt_rsc_1_4_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_4_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_4_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_4_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_4_i_1_inst_xt_rsc_1_4_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_4_i_1_inst_xt_rsc_1_4_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_5_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_5_i_oswt : IN STD_LOGIC;
      xt_rsc_1_5_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_5_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_5_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_5_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_5_i_1_inst_xt_rsc_1_5_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_5_i_1_inst_xt_rsc_1_5_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_6_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_6_i_oswt : IN STD_LOGIC;
      xt_rsc_1_6_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_6_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_6_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_6_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_6_i_1_inst_xt_rsc_1_6_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_6_i_1_inst_xt_rsc_1_6_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_7_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_7_i_oswt : IN STD_LOGIC;
      xt_rsc_1_7_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_7_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_7_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_7_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_7_i_1_inst_xt_rsc_1_7_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_7_i_1_inst_xt_rsc_1_7_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_8_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_8_i_oswt : IN STD_LOGIC;
      xt_rsc_1_8_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_8_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_8_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_8_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_8_i_1_inst_xt_rsc_1_8_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_8_i_1_inst_xt_rsc_1_8_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_9_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_9_i_oswt : IN STD_LOGIC;
      xt_rsc_1_9_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_9_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_9_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_9_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_9_i_1_inst_xt_rsc_1_9_i_qa_d : STD_LOGIC_VECTOR (31
      DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_9_i_1_inst_xt_rsc_1_9_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_10_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_10_i_oswt : IN STD_LOGIC;
      xt_rsc_1_10_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_10_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_10_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_10_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_10_i_1_inst_xt_rsc_1_10_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_10_i_1_inst_xt_rsc_1_10_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_11_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_11_i_oswt : IN STD_LOGIC;
      xt_rsc_1_11_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_11_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_11_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_11_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_11_i_1_inst_xt_rsc_1_11_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_11_i_1_inst_xt_rsc_1_11_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_12_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_12_i_oswt : IN STD_LOGIC;
      xt_rsc_1_12_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_12_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_12_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_12_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_12_i_1_inst_xt_rsc_1_12_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_12_i_1_inst_xt_rsc_1_12_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_13_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_13_i_oswt : IN STD_LOGIC;
      xt_rsc_1_13_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_13_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_13_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_13_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_13_i_1_inst_xt_rsc_1_13_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_13_i_1_inst_xt_rsc_1_13_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_14_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_14_i_oswt : IN STD_LOGIC;
      xt_rsc_1_14_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_14_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_14_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_14_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_14_i_1_inst_xt_rsc_1_14_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_14_i_1_inst_xt_rsc_1_14_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_15_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_15_i_oswt : IN STD_LOGIC;
      xt_rsc_1_15_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_15_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_15_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_15_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_15_i_1_inst_xt_rsc_1_15_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_15_i_1_inst_xt_rsc_1_15_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_16_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_16_i_oswt : IN STD_LOGIC;
      xt_rsc_1_16_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_16_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_16_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_16_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_16_i_1_inst_xt_rsc_1_16_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_16_i_1_inst_xt_rsc_1_16_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_17_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_17_i_oswt : IN STD_LOGIC;
      xt_rsc_1_17_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_17_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_17_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_17_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_17_i_1_inst_xt_rsc_1_17_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_17_i_1_inst_xt_rsc_1_17_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_18_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_18_i_oswt : IN STD_LOGIC;
      xt_rsc_1_18_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_18_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_18_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_18_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_18_i_1_inst_xt_rsc_1_18_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_18_i_1_inst_xt_rsc_1_18_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_19_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_19_i_oswt : IN STD_LOGIC;
      xt_rsc_1_19_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_19_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_19_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_19_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_19_i_1_inst_xt_rsc_1_19_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_19_i_1_inst_xt_rsc_1_19_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_20_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_20_i_oswt : IN STD_LOGIC;
      xt_rsc_1_20_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_20_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_20_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_20_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_20_i_1_inst_xt_rsc_1_20_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_20_i_1_inst_xt_rsc_1_20_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_21_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_21_i_oswt : IN STD_LOGIC;
      xt_rsc_1_21_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_21_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_21_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_21_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_21_i_1_inst_xt_rsc_1_21_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_21_i_1_inst_xt_rsc_1_21_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_22_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_22_i_oswt : IN STD_LOGIC;
      xt_rsc_1_22_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_22_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_22_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_22_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_22_i_1_inst_xt_rsc_1_22_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_22_i_1_inst_xt_rsc_1_22_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_23_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_23_i_oswt : IN STD_LOGIC;
      xt_rsc_1_23_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_23_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_23_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_23_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_23_i_1_inst_xt_rsc_1_23_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_23_i_1_inst_xt_rsc_1_23_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_24_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_24_i_oswt : IN STD_LOGIC;
      xt_rsc_1_24_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_24_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_24_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_24_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_24_i_1_inst_xt_rsc_1_24_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_24_i_1_inst_xt_rsc_1_24_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_25_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_25_i_oswt : IN STD_LOGIC;
      xt_rsc_1_25_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_25_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_25_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_25_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_25_i_1_inst_xt_rsc_1_25_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_25_i_1_inst_xt_rsc_1_25_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_26_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_26_i_oswt : IN STD_LOGIC;
      xt_rsc_1_26_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_26_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_26_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_26_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_26_i_1_inst_xt_rsc_1_26_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_26_i_1_inst_xt_rsc_1_26_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_27_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_27_i_oswt : IN STD_LOGIC;
      xt_rsc_1_27_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_27_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_27_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_27_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_27_i_1_inst_xt_rsc_1_27_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_27_i_1_inst_xt_rsc_1_27_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_28_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_28_i_oswt : IN STD_LOGIC;
      xt_rsc_1_28_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_28_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_28_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_28_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_28_i_1_inst_xt_rsc_1_28_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_28_i_1_inst_xt_rsc_1_28_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_29_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_29_i_oswt : IN STD_LOGIC;
      xt_rsc_1_29_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_29_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_29_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_29_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_29_i_1_inst_xt_rsc_1_29_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_29_i_1_inst_xt_rsc_1_29_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_30_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_30_i_oswt : IN STD_LOGIC;
      xt_rsc_1_30_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_30_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_30_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_30_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_30_i_1_inst_xt_rsc_1_30_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_30_i_1_inst_xt_rsc_1_30_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_1_31_i_1
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_1_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      core_wen : IN STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_1_31_i_oswt : IN STD_LOGIC;
      xt_rsc_1_31_i_qa_d_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct : IN STD_LOGIC;
      xt_rsc_1_31_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_31_i_wea_d_core_psct_pff : IN STD_LOGIC;
      xt_rsc_1_31_i_oswt_pff : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_xt_rsc_1_31_i_1_inst_xt_rsc_1_31_i_qa_d : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_xt_rsc_1_31_i_1_inst_xt_rsc_1_31_i_qa_d_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_0_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_0_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_0_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_0_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_0_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_0_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_0_RID : OUT STD_LOGIC;
      twiddle_rsc_0_0_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_0_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_0_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_0_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_0_ARID : IN STD_LOGIC;
      twiddle_rsc_0_0_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_0_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_0_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_0_BID : OUT STD_LOGIC;
      twiddle_rsc_0_0_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_0_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_0_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_0_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_0_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_0_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_0_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_0_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_0_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_0_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_i_s_raddr_core : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_1_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_1_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_1_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_1_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_1_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_1_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_1_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_1_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_1_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_1_RID : OUT STD_LOGIC;
      twiddle_rsc_0_1_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_1_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_1_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_1_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_1_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_1_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_1_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_1_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_1_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_1_ARID : IN STD_LOGIC;
      twiddle_rsc_0_1_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_1_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_1_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_1_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_1_BID : OUT STD_LOGIC;
      twiddle_rsc_0_1_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_1_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_1_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_1_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_1_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_1_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_1_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_1_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_1_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_1_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_1_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_1_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_1_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_1_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_1_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_1_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_1_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_1_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_1_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_i_s_raddr_core : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_2_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_2_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_2_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_2_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_2_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_2_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_2_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_2_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_2_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_2_RID : OUT STD_LOGIC;
      twiddle_rsc_0_2_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_2_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_2_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_2_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_2_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_2_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_2_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_2_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_2_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_2_ARID : IN STD_LOGIC;
      twiddle_rsc_0_2_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_2_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_2_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_2_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_2_BID : OUT STD_LOGIC;
      twiddle_rsc_0_2_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_2_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_2_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_2_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_2_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_2_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_2_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_2_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_2_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_2_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_2_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_2_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_2_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_2_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_2_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_2_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_2_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_2_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_2_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_i_s_raddr_core : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_3_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_3_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_3_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_3_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_3_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_3_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_3_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_3_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_3_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_3_RID : OUT STD_LOGIC;
      twiddle_rsc_0_3_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_3_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_3_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_3_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_3_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_3_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_3_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_3_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_3_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_3_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_3_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_3_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_3_ARID : IN STD_LOGIC;
      twiddle_rsc_0_3_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_3_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_3_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_3_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_3_BID : OUT STD_LOGIC;
      twiddle_rsc_0_3_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_3_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_3_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_3_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_3_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_3_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_3_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_3_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_3_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_3_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_3_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_3_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_3_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_3_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_3_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_3_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_3_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_3_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_3_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_3_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_3_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_3_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_3_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_i_s_raddr_core : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_4_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_4_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_4_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_4_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_4_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_4_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_4_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_4_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_4_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_4_RID : OUT STD_LOGIC;
      twiddle_rsc_0_4_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_4_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_4_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_4_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_4_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_4_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_4_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_4_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_4_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_4_ARID : IN STD_LOGIC;
      twiddle_rsc_0_4_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_4_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_4_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_4_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_4_BID : OUT STD_LOGIC;
      twiddle_rsc_0_4_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_4_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_4_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_4_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_4_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_4_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_4_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_4_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_4_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_4_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_4_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_4_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_4_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_4_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_4_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_4_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_4_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_4_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_4_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_i_s_raddr_core : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_5_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_5_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_5_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_5_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_5_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_5_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_5_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_5_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_5_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_5_RID : OUT STD_LOGIC;
      twiddle_rsc_0_5_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_5_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_5_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_5_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_5_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_5_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_5_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_5_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_5_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_5_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_5_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_5_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_5_ARID : IN STD_LOGIC;
      twiddle_rsc_0_5_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_5_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_5_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_5_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_5_BID : OUT STD_LOGIC;
      twiddle_rsc_0_5_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_5_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_5_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_5_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_5_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_5_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_5_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_5_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_5_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_5_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_5_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_5_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_5_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_5_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_5_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_5_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_5_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_5_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_5_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_5_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_5_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_5_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_5_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_i_s_raddr_core : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_6_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_6_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_6_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_6_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_6_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_6_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_6_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_6_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_6_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_6_RID : OUT STD_LOGIC;
      twiddle_rsc_0_6_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_6_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_6_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_6_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_6_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_6_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_6_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_6_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_6_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_6_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_6_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_6_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_6_ARID : IN STD_LOGIC;
      twiddle_rsc_0_6_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_6_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_6_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_6_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_6_BID : OUT STD_LOGIC;
      twiddle_rsc_0_6_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_6_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_6_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_6_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_6_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_6_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_6_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_6_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_6_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_6_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_6_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_6_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_6_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_6_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_6_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_6_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_6_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_6_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_6_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_6_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_6_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_6_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_6_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_i_s_raddr_core : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_7_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_7_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_7_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_7_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_7_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_7_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_7_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_7_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_7_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_7_RID : OUT STD_LOGIC;
      twiddle_rsc_0_7_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_7_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_7_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_7_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_7_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_7_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_7_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_7_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_7_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_7_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_7_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_7_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_7_ARID : IN STD_LOGIC;
      twiddle_rsc_0_7_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_7_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_7_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_7_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_7_BID : OUT STD_LOGIC;
      twiddle_rsc_0_7_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_7_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_7_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_7_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_7_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_7_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_7_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_7_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_7_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_7_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_7_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_7_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_7_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_7_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_7_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_7_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_7_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_7_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_7_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_7_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_7_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_7_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_7_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_i_s_raddr_core : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_8_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_8_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_8_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_8_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_8_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_8_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_8_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_8_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_8_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_8_RID : OUT STD_LOGIC;
      twiddle_rsc_0_8_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_8_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_8_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_8_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_8_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_8_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_8_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_8_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_8_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_8_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_8_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_8_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_8_ARID : IN STD_LOGIC;
      twiddle_rsc_0_8_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_8_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_8_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_8_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_8_BID : OUT STD_LOGIC;
      twiddle_rsc_0_8_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_8_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_8_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_8_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_8_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_8_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_8_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_8_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_8_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_8_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_8_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_8_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_8_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_8_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_8_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_8_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_8_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_8_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_8_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_8_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_8_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_8_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_8_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_i_s_raddr_core : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_9_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_9_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_9_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_9_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_9_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_9_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_9_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_9_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_9_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_9_RID : OUT STD_LOGIC;
      twiddle_rsc_0_9_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_9_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_9_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_9_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_9_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_9_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_9_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_9_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_9_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_9_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_9_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_9_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_9_ARID : IN STD_LOGIC;
      twiddle_rsc_0_9_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_9_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_9_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_9_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_9_BID : OUT STD_LOGIC;
      twiddle_rsc_0_9_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_9_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_9_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_9_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_9_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_9_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_9_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_9_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_9_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_9_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_9_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_9_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_9_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_9_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_9_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_9_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_9_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_9_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_9_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_9_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_9_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_9_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_9_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_i_s_raddr_core : STD_LOGIC_VECTOR
      (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_10_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_10_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_10_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_10_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_10_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_10_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_10_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_10_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_10_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_10_RID : OUT STD_LOGIC;
      twiddle_rsc_0_10_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_10_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_10_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_10_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_10_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_10_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_10_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_10_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_10_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_10_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_10_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_10_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_10_ARID : IN STD_LOGIC;
      twiddle_rsc_0_10_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_10_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_10_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_10_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_10_BID : OUT STD_LOGIC;
      twiddle_rsc_0_10_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_10_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_10_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_10_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_10_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_10_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_10_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_10_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_10_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_10_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_10_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_10_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_10_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_10_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_10_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_10_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_10_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_10_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_10_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_10_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_10_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_10_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_10_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_i_s_raddr_core :
      STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_11_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_11_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_11_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_11_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_11_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_11_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_11_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_11_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_11_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_11_RID : OUT STD_LOGIC;
      twiddle_rsc_0_11_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_11_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_11_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_11_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_11_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_11_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_11_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_11_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_11_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_11_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_11_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_11_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_11_ARID : IN STD_LOGIC;
      twiddle_rsc_0_11_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_11_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_11_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_11_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_11_BID : OUT STD_LOGIC;
      twiddle_rsc_0_11_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_11_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_11_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_11_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_11_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_11_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_11_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_11_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_11_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_11_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_11_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_11_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_11_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_11_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_11_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_11_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_11_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_11_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_11_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_11_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_11_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_11_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_11_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_i_s_raddr_core :
      STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_12_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_12_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_12_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_12_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_12_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_12_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_12_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_12_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_12_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_12_RID : OUT STD_LOGIC;
      twiddle_rsc_0_12_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_12_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_12_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_12_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_12_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_12_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_12_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_12_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_12_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_12_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_12_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_12_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_12_ARID : IN STD_LOGIC;
      twiddle_rsc_0_12_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_12_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_12_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_12_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_12_BID : OUT STD_LOGIC;
      twiddle_rsc_0_12_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_12_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_12_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_12_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_12_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_12_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_12_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_12_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_12_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_12_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_12_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_12_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_12_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_12_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_12_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_12_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_12_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_12_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_12_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_12_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_12_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_12_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_12_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_i_s_raddr_core :
      STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_13_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_13_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_13_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_13_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_13_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_13_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_13_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_13_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_13_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_13_RID : OUT STD_LOGIC;
      twiddle_rsc_0_13_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_13_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_13_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_13_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_13_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_13_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_13_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_13_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_13_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_13_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_13_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_13_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_13_ARID : IN STD_LOGIC;
      twiddle_rsc_0_13_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_13_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_13_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_13_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_13_BID : OUT STD_LOGIC;
      twiddle_rsc_0_13_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_13_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_13_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_13_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_13_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_13_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_13_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_13_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_13_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_13_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_13_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_13_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_13_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_13_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_13_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_13_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_13_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_13_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_13_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_13_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_13_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_13_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_13_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_i_s_raddr_core :
      STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_14_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_14_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_14_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_14_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_14_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_14_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_14_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_14_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_14_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_14_RID : OUT STD_LOGIC;
      twiddle_rsc_0_14_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_14_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_14_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_14_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_14_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_14_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_14_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_14_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_14_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_14_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_14_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_14_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_14_ARID : IN STD_LOGIC;
      twiddle_rsc_0_14_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_14_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_14_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_14_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_14_BID : OUT STD_LOGIC;
      twiddle_rsc_0_14_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_14_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_14_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_14_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_14_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_14_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_14_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_14_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_14_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_14_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_14_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_14_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_14_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_14_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_14_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_14_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_14_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_14_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_14_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_14_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_14_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_14_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_14_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_i_s_raddr_core :
      STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_rsc_0_15_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_rsc_0_15_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_15_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_15_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_15_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_15_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_15_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_15_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_15_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_15_RID : OUT STD_LOGIC;
      twiddle_rsc_0_15_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_15_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_15_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_15_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_15_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_15_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_15_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_15_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_15_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_15_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_15_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_15_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_15_ARID : IN STD_LOGIC;
      twiddle_rsc_0_15_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_15_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_15_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_15_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_15_BID : OUT STD_LOGIC;
      twiddle_rsc_0_15_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_15_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_15_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_15_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_15_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_15_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_15_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_15_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_15_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_15_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_15_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_15_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_15_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_15_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_15_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_15_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_15_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_15_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_15_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_rsc_0_15_i_oswt : IN STD_LOGIC;
      twiddle_rsc_0_15_i_wen_comp : OUT STD_LOGIC;
      twiddle_rsc_0_15_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_rsc_0_15_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_i_s_raddr_core :
      STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_i_s_din_mxwt : STD_LOGIC_VECTOR
      (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_0_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_0_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_0_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_0_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_0_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_0_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_0_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_0_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_0_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_0_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_0_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_0_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_0_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_0_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_0_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_0_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_0_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_0_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_0_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_1_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_1_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_1_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_1_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_1_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_1_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_1_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_1_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_1_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_1_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_1_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_1_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_1_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_1_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_1_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_1_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_1_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_1_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_1_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_1_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_1_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_1_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_1_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_1_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_1_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_1_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_1_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_1_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_1_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_1_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_1_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_1_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_1_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_1_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_1_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_1_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_1_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_1_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_2_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_2_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_2_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_2_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_2_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_2_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_2_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_2_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_2_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_2_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_2_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_2_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_2_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_2_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_2_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_2_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_2_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_2_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_2_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_2_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_2_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_2_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_2_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_2_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_2_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_2_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_2_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_2_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_2_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_2_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_2_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_2_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_2_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_2_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_2_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_2_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_2_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_2_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_3_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_3_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_3_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_3_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_3_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_3_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_3_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_3_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_3_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_3_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_3_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_3_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_3_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_3_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_3_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_3_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_3_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_3_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_3_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_3_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_3_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_3_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_3_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_3_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_3_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_3_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_3_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_3_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_3_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_3_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_3_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_3_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_3_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_3_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_3_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_3_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_3_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_3_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_4_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_4_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_4_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_4_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_4_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_4_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_4_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_4_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_4_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_4_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_4_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_4_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_4_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_4_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_4_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_4_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_4_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_4_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_4_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_4_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_4_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_4_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_4_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_4_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_4_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_4_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_4_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_4_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_4_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_4_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_4_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_4_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_4_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_4_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_4_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_4_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_4_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_4_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_5_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_5_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_5_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_5_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_5_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_5_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_5_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_5_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_5_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_5_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_5_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_5_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_5_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_5_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_5_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_5_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_5_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_5_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_5_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_5_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_5_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_5_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_5_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_5_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_5_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_5_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_5_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_5_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_5_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_5_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_5_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_5_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_5_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_5_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_5_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_5_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_5_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_5_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_6_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_6_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_6_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_6_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_6_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_6_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_6_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_6_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_6_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_6_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_6_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_6_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_6_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_6_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_6_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_6_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_6_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_6_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_6_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_6_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_6_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_6_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_6_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_6_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_6_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_6_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_6_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_6_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_6_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_6_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_6_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_6_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_6_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_6_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_6_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_6_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_6_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_6_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_7_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_7_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_7_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_7_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_7_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_7_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_7_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_7_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_7_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_7_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_7_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_7_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_7_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_7_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_7_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_7_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_7_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_7_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_7_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_7_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_7_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_7_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_7_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_7_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_7_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_7_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_7_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_7_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_7_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_7_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_7_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_7_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_7_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_7_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_7_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_7_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_7_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_7_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_8_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_8_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_8_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_8_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_8_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_8_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_8_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_8_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_8_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_8_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_8_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_8_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_8_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_8_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_8_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_8_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_8_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_8_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_8_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_8_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_8_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_8_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_8_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_8_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_8_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_8_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_8_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_8_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_8_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_8_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_8_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_8_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_8_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_8_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_8_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_8_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_8_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_8_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_8_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_8_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_9_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_9_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_9_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_9_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_9_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_9_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_9_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_9_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_9_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_9_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_9_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_9_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_9_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_9_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_9_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_9_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_9_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_9_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_9_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_9_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_9_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_9_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_9_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_9_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_9_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_9_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_9_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_9_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_9_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_9_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_9_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_9_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_9_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_9_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_9_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_9_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_9_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_9_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_9_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_9_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_i_s_din_mxwt :
      STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_10_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_10_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_10_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_10_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_10_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_10_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_10_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_10_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_10_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_10_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_10_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_10_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_10_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_10_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_10_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_10_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_10_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_10_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_10_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_10_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_10_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_10_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_10_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_10_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_10_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_10_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_10_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_10_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_10_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_10_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_10_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_10_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_10_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_10_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_10_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_10_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_10_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_10_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_10_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_10_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_11_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_11_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_11_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_11_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_11_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_11_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_11_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_11_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_11_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_11_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_11_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_11_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_11_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_11_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_11_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_11_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_11_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_11_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_11_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_11_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_11_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_11_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_11_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_11_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_11_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_11_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_11_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_11_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_11_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_11_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_11_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_11_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_11_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_11_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_11_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_11_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_11_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_11_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_11_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_11_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_12_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_12_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_12_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_12_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_12_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_12_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_12_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_12_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_12_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_12_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_12_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_12_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_12_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_12_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_12_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_12_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_12_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_12_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_12_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_12_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_12_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_12_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_12_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_12_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_12_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_12_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_12_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_12_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_12_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_12_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_12_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_12_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_12_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_12_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_12_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_12_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_12_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_12_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_12_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_12_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_13_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_13_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_13_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_13_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_13_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_13_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_13_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_13_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_13_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_13_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_13_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_13_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_13_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_13_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_13_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_13_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_13_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_13_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_13_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_13_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_13_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_13_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_13_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_13_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_13_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_13_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_13_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_13_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_13_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_13_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_13_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_13_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_13_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_13_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_13_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_13_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_13_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_13_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_13_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_13_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_14_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_14_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_14_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_14_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_14_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_14_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_14_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_14_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_14_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_14_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_14_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_14_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_14_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_14_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_14_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_14_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_14_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_14_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_14_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_14_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_14_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_14_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_14_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_14_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_14_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_14_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_14_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_14_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_14_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_14_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_14_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_14_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_14_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_14_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_14_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_14_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_14_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_14_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_14_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_14_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_twiddle_h_rsc_0_15_i
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      twiddle_h_rsc_0_15_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_15_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_15_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_15_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_15_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_15_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_15_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_15_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_15_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_15_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_15_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_15_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_15_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_15_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_15_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_15_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_15_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_15_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_15_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_15_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_15_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_15_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_15_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_15_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_15_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_15_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_15_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_15_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_15_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_15_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_15_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_15_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_15_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_15_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_15_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_15_AWID : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      twiddle_h_rsc_0_15_i_oswt : IN STD_LOGIC;
      twiddle_h_rsc_0_15_i_wen_comp : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_i_s_raddr_core : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
      twiddle_h_rsc_0_15_i_s_din_mxwt : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_RRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_RDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_BRESP : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_WSTRB : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_WDATA : STD_LOGIC_VECTOR
      (31 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWREGION : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWQOS : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWPROT : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWCACHE : STD_LOGIC_VECTOR
      (3 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWBURST : STD_LOGIC_VECTOR
      (1 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWSIZE : STD_LOGIC_VECTOR
      (2 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWLEN : STD_LOGIC_VECTOR
      (7 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWADDR : STD_LOGIC_VECTOR
      (11 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_i_s_raddr_core
      : STD_LOGIC_VECTOR (5 DOWNTO 0);
  SIGNAL peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_i_s_din_mxwt
      : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core_xt_rsc_triosy_1_31_obj
    PORT(
      xt_rsc_triosy_1_31_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_31_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_30_obj
    PORT(
      xt_rsc_triosy_1_30_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_30_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_29_obj
    PORT(
      xt_rsc_triosy_1_29_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_29_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_28_obj
    PORT(
      xt_rsc_triosy_1_28_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_28_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_27_obj
    PORT(
      xt_rsc_triosy_1_27_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_27_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_26_obj
    PORT(
      xt_rsc_triosy_1_26_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_26_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_25_obj
    PORT(
      xt_rsc_triosy_1_25_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_25_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_24_obj
    PORT(
      xt_rsc_triosy_1_24_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_24_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_23_obj
    PORT(
      xt_rsc_triosy_1_23_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_23_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_22_obj
    PORT(
      xt_rsc_triosy_1_22_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_22_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_21_obj
    PORT(
      xt_rsc_triosy_1_21_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_21_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_20_obj
    PORT(
      xt_rsc_triosy_1_20_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_20_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_19_obj
    PORT(
      xt_rsc_triosy_1_19_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_19_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_18_obj
    PORT(
      xt_rsc_triosy_1_18_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_18_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_17_obj
    PORT(
      xt_rsc_triosy_1_17_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_17_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_16_obj
    PORT(
      xt_rsc_triosy_1_16_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_16_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_15_obj
    PORT(
      xt_rsc_triosy_1_15_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_15_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_14_obj
    PORT(
      xt_rsc_triosy_1_14_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_14_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_13_obj
    PORT(
      xt_rsc_triosy_1_13_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_13_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_12_obj
    PORT(
      xt_rsc_triosy_1_12_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_12_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_11_obj
    PORT(
      xt_rsc_triosy_1_11_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_11_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_10_obj
    PORT(
      xt_rsc_triosy_1_10_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_10_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_9_obj
    PORT(
      xt_rsc_triosy_1_9_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_9_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_8_obj
    PORT(
      xt_rsc_triosy_1_8_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_8_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_7_obj
    PORT(
      xt_rsc_triosy_1_7_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_7_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_6_obj
    PORT(
      xt_rsc_triosy_1_6_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_6_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_5_obj
    PORT(
      xt_rsc_triosy_1_5_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_5_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_4_obj
    PORT(
      xt_rsc_triosy_1_4_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_4_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_3_obj
    PORT(
      xt_rsc_triosy_1_3_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_3_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_2_obj
    PORT(
      xt_rsc_triosy_1_2_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_2_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_1_obj
    PORT(
      xt_rsc_triosy_1_1_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_1_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_1_0_obj
    PORT(
      xt_rsc_triosy_1_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_1_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_31_obj
    PORT(
      xt_rsc_triosy_0_31_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_31_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_30_obj
    PORT(
      xt_rsc_triosy_0_30_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_30_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_29_obj
    PORT(
      xt_rsc_triosy_0_29_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_29_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_28_obj
    PORT(
      xt_rsc_triosy_0_28_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_28_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_27_obj
    PORT(
      xt_rsc_triosy_0_27_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_27_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_26_obj
    PORT(
      xt_rsc_triosy_0_26_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_26_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_25_obj
    PORT(
      xt_rsc_triosy_0_25_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_25_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_24_obj
    PORT(
      xt_rsc_triosy_0_24_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_24_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_23_obj
    PORT(
      xt_rsc_triosy_0_23_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_23_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_22_obj
    PORT(
      xt_rsc_triosy_0_22_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_22_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_21_obj
    PORT(
      xt_rsc_triosy_0_21_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_21_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_20_obj
    PORT(
      xt_rsc_triosy_0_20_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_20_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_19_obj
    PORT(
      xt_rsc_triosy_0_19_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_19_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_18_obj
    PORT(
      xt_rsc_triosy_0_18_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_18_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_17_obj
    PORT(
      xt_rsc_triosy_0_17_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_17_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_16_obj
    PORT(
      xt_rsc_triosy_0_16_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_16_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_15_obj
    PORT(
      xt_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_15_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_14_obj
    PORT(
      xt_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_14_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_13_obj
    PORT(
      xt_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_13_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_12_obj
    PORT(
      xt_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_12_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_11_obj
    PORT(
      xt_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_11_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_10_obj
    PORT(
      xt_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_10_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_9_obj
    PORT(
      xt_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_9_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_8_obj
    PORT(
      xt_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_8_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_7_obj
    PORT(
      xt_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_6_obj
    PORT(
      xt_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_5_obj
    PORT(
      xt_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_4_obj
    PORT(
      xt_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_3_obj
    PORT(
      xt_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_2_obj
    PORT(
      xt_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_1_obj
    PORT(
      xt_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_xt_rsc_triosy_0_0_obj
    PORT(
      xt_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      xt_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_p_rsc_triosy_obj
    PORT(
      p_rsc_triosy_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      p_rsc_triosy_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_r_rsc_triosy_obj
    PORT(
      r_rsc_triosy_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      r_rsc_triosy_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_15_obj
    PORT(
      twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_15_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_14_obj
    PORT(
      twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_14_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_13_obj
    PORT(
      twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_13_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_12_obj
    PORT(
      twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_12_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_11_obj
    PORT(
      twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_11_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_10_obj
    PORT(
      twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_10_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_9_obj
    PORT(
      twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_9_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_8_obj
    PORT(
      twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_8_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_7_obj
    PORT(
      twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_6_obj
    PORT(
      twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_5_obj
    PORT(
      twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_4_obj
    PORT(
      twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_3_obj
    PORT(
      twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_2_obj
    PORT(
      twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_1_obj
    PORT(
      twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_rsc_triosy_0_0_obj
    PORT(
      twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_15_obj
    PORT(
      twiddle_h_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_15_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_14_obj
    PORT(
      twiddle_h_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_14_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_13_obj
    PORT(
      twiddle_h_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_13_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_12_obj
    PORT(
      twiddle_h_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_12_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_11_obj
    PORT(
      twiddle_h_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_11_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_10_obj
    PORT(
      twiddle_h_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_10_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_9_obj
    PORT(
      twiddle_h_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_9_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_8_obj
    PORT(
      twiddle_h_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_8_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_7_obj
    PORT(
      twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_7_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_6_obj
    PORT(
      twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_6_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_5_obj
    PORT(
      twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_5_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_4_obj
    PORT(
      twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_4_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_3_obj
    PORT(
      twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_3_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_2_obj
    PORT(
      twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_2_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_1_obj
    PORT(
      twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_1_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_twiddle_h_rsc_triosy_0_0_obj
    PORT(
      twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      core_wten : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_0_obj_iswt0 : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_staller
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      core_wen : OUT STD_LOGIC;
      core_wten : OUT STD_LOGIC;
      twiddle_rsc_0_0_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_1_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_2_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_3_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_4_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_5_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_6_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_7_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_8_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_9_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_10_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_11_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_12_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_13_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_14_i_wen_comp : IN STD_LOGIC;
      twiddle_rsc_0_15_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_0_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_1_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_2_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_3_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_4_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_5_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_6_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_7_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_8_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_9_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_10_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_11_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_12_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_13_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_14_i_wen_comp : IN STD_LOGIC;
      twiddle_h_rsc_0_15_i_wen_comp : IN STD_LOGIC
    );
  END COMPONENT;
  COMPONENT peaseNTT_core_core_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      core_wen : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (9 DOWNTO 0);
      INNER_LOOP1_C_0_tr0 : IN STD_LOGIC;
      INNER_LOOP2_C_0_tr0 : IN STD_LOGIC;
      INNER_LOOP2_C_0_tr1 : IN STD_LOGIC;
      INNER_LOOP3_C_0_tr0 : IN STD_LOGIC;
      INNER_LOOP4_C_0_tr0 : IN STD_LOGIC;
      INNER_LOOP4_C_0_tr1 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_core_fsm_inst_fsm_output : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL peaseNTT_core_core_fsm_inst_INNER_LOOP2_C_0_tr0 : STD_LOGIC;
  SIGNAL peaseNTT_core_core_fsm_inst_INNER_LOOP2_C_0_tr1 : STD_LOGIC;
  SIGNAL peaseNTT_core_core_fsm_inst_INNER_LOOP3_C_0_tr0 : STD_LOGIC;
  SIGNAL peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX1HOT_s_1_4_2(input_3 : STD_LOGIC;
  input_2 : STD_LOGIC;
  input_1 : STD_LOGIC;
  input_0 : STD_LOGIC;
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;
    VARIABLE tmp : STD_LOGIC;

    BEGIN
      tmp := sel(0);
      result := input_0 and tmp;
      tmp := sel(1);
      result := result or ( input_1 and tmp);
      tmp := sel(2);
      result := result or ( input_2 and tmp);
      tmp := sel(3);
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_2_4_2(input_3 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(1 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(1 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(1 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_31_4_2(input_3 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(30 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(30 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_12_2(input_11 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_10 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_9 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(11 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
      tmp := (OTHERS=>sel( 9));
      result := result or ( input_9 and tmp);
      tmp := (OTHERS=>sel( 10));
      result := result or ( input_10 and tmp);
      tmp := (OTHERS=>sel( 11));
      result := result or ( input_11 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_3_2(input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_4_2(input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_5_2(input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(4 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_6_2(input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(5 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_8_2(input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(7 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_32_9_2(input_8 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_7 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_6 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_5 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_4 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(8 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
      tmp := (OTHERS=>sel( 4));
      result := result or ( input_4 and tmp);
      tmp := (OTHERS=>sel( 5));
      result := result or ( input_5 and tmp);
      tmp := (OTHERS=>sel( 6));
      result := result or ( input_6 and tmp);
      tmp := (OTHERS=>sel( 7));
      result := result or ( input_7 and tmp);
      tmp := (OTHERS=>sel( 8));
      result := result or ( input_8 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_3_3_2(input_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(2 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
    RETURN result;
  END;

  FUNCTION MUX1HOT_v_4_4_2(input_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC_VECTOR(3 DOWNTO 0))
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE tmp : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      tmp := (OTHERS=>sel(0));
      result := input_0 and tmp;
      tmp := (OTHERS=>sel( 1));
      result := result or ( input_1 and tmp);
      tmp := (OTHERS=>sel( 2));
      result := result or ( input_2 and tmp);
      tmp := (OTHERS=>sel( 3));
      result := result or ( input_3 and tmp);
    RETURN result;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_31_2_2(input_0 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(30 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(30 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_32_2_2(input_0 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(31 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_5_2_2(input_0 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(4 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(4 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

BEGIN
  p_rsci : work.ccs_in_pkg_v1.ccs_in_v1
    GENERIC MAP(
      rscid => 2,
      width => 32
      )
    PORT MAP(
      dat => p_rsci_dat,
      idat => p_rsci_idat_1
    );
  p_rsci_dat <= p_rsc_dat;
  p_rsci_idat <= p_rsci_idat_1;

  mult_t_mul_cmp : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_a,
      b => mult_t_mul_cmp_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_z_1
    );
  mult_t_mul_cmp_a <= MUX1HOT_v_32_4_2(tmp_65_lpi_3_dfm_mx0, tmp_1_lpi_3_dfm_mx0,
      mult_t_mul_cmp_a_mx0w2, tmp_31_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_b <= MUX1HOT_v_32_9_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_8_i_s_din_mxwt,
      twiddle_h_rsc_0_9_i_s_din_mxwt, twiddle_h_rsc_0_10_i_s_din_mxwt, twiddle_h_rsc_0_11_i_s_din_mxwt,
      twiddle_h_rsc_0_12_i_s_din_mxwt, twiddle_h_rsc_0_13_i_s_din_mxwt, twiddle_h_rsc_0_14_i_s_din_mxwt,
      twiddle_h_rsc_0_15_i_s_din_mxwt, STD_LOGIC_VECTOR'( or_dcpl_29 & INNER_LOOP1_tw_h_and_44_cse
      & INNER_LOOP1_tw_h_and_45_cse & INNER_LOOP1_tw_h_and_46_cse & INNER_LOOP1_tw_h_and_47_cse
      & INNER_LOOP1_tw_h_or_9_cse & INNER_LOOP1_tw_h_or_10_cse & INNER_LOOP1_tw_h_or_11_cse
      & INNER_LOOP1_tw_h_or_12_cse));
  mult_t_mul_cmp_z <= mult_t_mul_cmp_z_1;

  mult_t_mul_cmp_1 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_1_a,
      b => mult_t_mul_cmp_1_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_1_z_1
    );
  mult_t_mul_cmp_1_a <= MUX1HOT_v_32_4_2(mult_t_mul_cmp_1_a_mx0w0, tmp_31_lpi_3_dfm_mx0,
      tmp_125_lpi_3_dfm_mx0, tmp_1_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_1_b <= MUX1HOT_v_32_5_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_8_i_s_din_mxwt,
      twiddle_h_rsc_0_10_i_s_din_mxwt, twiddle_h_rsc_0_12_i_s_din_mxwt, twiddle_h_rsc_0_14_i_s_din_mxwt,
      STD_LOGIC_VECTOR'( (NOT (fsm_output(6))) & INNER_LOOP1_tw_h_and_40_cse & INNER_LOOP1_tw_h_and_41_cse
      & INNER_LOOP1_tw_h_and_42_cse & INNER_LOOP1_tw_h_and_43_cse));
  mult_t_mul_cmp_1_z <= mult_t_mul_cmp_1_z_1;

  mult_t_mul_cmp_2 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_2_a,
      b => mult_t_mul_cmp_2_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_2_z_1
    );
  mult_t_mul_cmp_2_a <= MUX1HOT_v_32_4_2(tmp_93_lpi_3_dfm_mx0, tmp_29_lpi_3_dfm_mx0,
      mult_t_mul_cmp_2_a_mx0w2, tmp_3_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_2_b <= MUX1HOT_v_32_6_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_8_i_s_din_mxwt,
      twiddle_h_rsc_0_9_i_s_din_mxwt, twiddle_h_rsc_0_12_i_s_din_mxwt, twiddle_h_rsc_0_13_i_s_din_mxwt,
      twiddle_h_rsc_0_1_i_s_din_mxwt, STD_LOGIC_VECTOR'( or_tmp_804 & INNER_LOOP1_tw_h_and_36_cse
      & INNER_LOOP1_tw_h_and_37_cse & INNER_LOOP1_tw_h_and_38_cse & INNER_LOOP1_tw_h_and_39_cse
      & or_tmp_806));
  mult_t_mul_cmp_2_z <= mult_t_mul_cmp_2_z_1;

  mult_t_mul_cmp_3 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_3_a,
      b => mult_t_mul_cmp_3_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_3_z_1
    );
  mult_t_mul_cmp_3_a <= MUX1HOT_v_32_4_2(tmp_91_lpi_3_dfm_mx0, tmp_27_lpi_3_dfm_mx0,
      tmp_121_lpi_3_dfm_mx0, tmp_5_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_3_b <= MUX1HOT_v_32_4_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_12_i_s_din_mxwt,
      twiddle_h_rsc_0_8_i_s_din_mxwt, twiddle_h_rsc_0_2_i_s_din_mxwt, STD_LOGIC_VECTOR'(
      (or_dcpl_29 OR and_1944_cse) & or_tmp_812 & and_1948_cse & or_tmp_814));
  mult_t_mul_cmp_3_z <= mult_t_mul_cmp_3_z_1;

  mult_t_mul_cmp_4 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_4_a,
      b => mult_t_mul_cmp_4_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_4_z_1
    );
  mult_t_mul_cmp_4_a <= MUX1HOT_v_32_4_2(tmp_89_lpi_3_dfm_mx0, tmp_25_lpi_3_dfm_mx0,
      mult_t_mul_cmp_4_a_mx0w2, tmp_7_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_4_b <= MUX1HOT_v_32_8_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_8_i_s_din_mxwt,
      twiddle_h_rsc_0_9_i_s_din_mxwt, twiddle_h_rsc_0_10_i_s_din_mxwt, twiddle_h_rsc_0_11_i_s_din_mxwt,
      twiddle_h_rsc_0_1_i_s_din_mxwt, twiddle_h_rsc_0_2_i_s_din_mxwt, twiddle_h_rsc_0_3_i_s_din_mxwt,
      STD_LOGIC_VECTOR'( (or_dcpl_29 OR INNER_LOOP1_tw_h_and_49_cse) & INNER_LOOP1_tw_h_and_29_cse
      & INNER_LOOP1_tw_h_and_30_cse & INNER_LOOP1_tw_h_and_31_cse & INNER_LOOP1_tw_h_and_32_cse
      & INNER_LOOP1_tw_h_and_51_cse & INNER_LOOP1_tw_h_and_53_cse & INNER_LOOP1_tw_h_and_55_cse));
  mult_t_mul_cmp_4_z <= mult_t_mul_cmp_4_z_1;

  mult_t_mul_cmp_5 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_5_a,
      b => mult_t_mul_cmp_5_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_5_z_1
    );
  mult_t_mul_cmp_5_a <= MUX1HOT_v_32_4_2(tmp_87_lpi_3_dfm_mx0, tmp_23_lpi_3_dfm_mx0,
      mult_t_mul_cmp_5_a_mx0w2, mult_t_mul_cmp_12_a_mx0w3, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_5_b <= MUX1HOT_v_32_4_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_10_i_s_din_mxwt,
      twiddle_h_rsc_0_8_i_s_din_mxwt, twiddle_h_rsc_0_4_i_s_din_mxwt, STD_LOGIC_VECTOR'(
      or_dcpl_29 & or_tmp_827 & and_1978_cse & (fsm_output(8))));
  mult_t_mul_cmp_5_z <= mult_t_mul_cmp_5_z_1;

  mult_t_mul_cmp_6 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_6_a,
      b => mult_t_mul_cmp_6_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_6_z_1
    );
  mult_t_mul_cmp_6_a <= MUX1HOT_v_32_4_2(tmp_85_lpi_3_dfm_mx0, tmp_21_lpi_3_dfm_mx0,
      mult_t_mul_cmp_6_a_mx0w2, mult_t_mul_cmp_11_a_mx0w3, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_6_b <= MUX1HOT_v_32_5_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_9_i_s_din_mxwt,
      twiddle_h_rsc_0_8_i_s_din_mxwt, twiddle_h_rsc_0_5_i_s_din_mxwt, twiddle_h_rsc_0_4_i_s_din_mxwt,
      STD_LOGIC_VECTOR'( or_dcpl_29 & or_tmp_835 & and_1994_cse & or_tmp_806 & and_1929_cse));
  mult_t_mul_cmp_6_z <= mult_t_mul_cmp_6_z_1;

  mult_t_mul_cmp_7 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_7_a,
      b => mult_t_mul_cmp_7_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_7_z_1
    );
  mult_t_mul_cmp_7_a <= MUX1HOT_v_32_4_2(tmp_83_lpi_3_dfm_mx0, tmp_19_lpi_3_dfm_mx0,
      mult_t_mul_cmp_7_a_mx0w2, mult_t_mul_cmp_10_a_mx0w3, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_7_b <= MUX1HOT_v_32_4_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_8_i_s_din_mxwt,
      twiddle_h_rsc_0_6_i_s_din_mxwt, twiddle_h_rsc_0_4_i_s_din_mxwt, STD_LOGIC_VECTOR'(
      or_dcpl_29 & (fsm_output(6)) & or_tmp_814 & and_1944_cse));
  mult_t_mul_cmp_7_z <= mult_t_mul_cmp_7_z_1;

  mult_t_mul_cmp_8 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_8_a,
      b => mult_t_mul_cmp_8_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_8_z_1
    );
  mult_t_mul_cmp_8_a <= MUX1HOT_v_32_4_2(tmp_81_lpi_3_dfm_mx0, tmp_17_lpi_3_dfm_mx0,
      mult_t_mul_cmp_8_a_mx0w2, mult_t_mul_cmp_9_a_mx0w3, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_8_b <= MUX1HOT_v_32_8_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_1_i_s_din_mxwt,
      twiddle_h_rsc_0_2_i_s_din_mxwt, twiddle_h_rsc_0_3_i_s_din_mxwt, twiddle_h_rsc_0_4_i_s_din_mxwt,
      twiddle_h_rsc_0_5_i_s_din_mxwt, twiddle_h_rsc_0_6_i_s_din_mxwt, twiddle_h_rsc_0_7_i_s_din_mxwt,
      STD_LOGIC_VECTOR'( INNER_LOOP1_tw_h_or_3_cse & INNER_LOOP1_tw_h_and_45_cse
      & INNER_LOOP1_tw_h_and_46_cse & INNER_LOOP1_tw_h_and_47_cse & INNER_LOOP1_tw_h_or_9_cse
      & INNER_LOOP1_tw_h_or_10_cse & INNER_LOOP1_tw_h_or_11_cse & INNER_LOOP1_tw_h_or_12_cse));
  mult_t_mul_cmp_8_z <= mult_t_mul_cmp_8_z_1;

  mult_t_mul_cmp_9 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_9_a,
      b => mult_t_mul_cmp_9_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_9_z_1
    );
  mult_t_mul_cmp_9_a <= MUX1HOT_v_32_4_2(mult_t_mul_cmp_9_a_mx0w0, mult_t_mul_cmp_9_a_mx0w3,
      mult_t_mul_cmp_9_a_mx0w2, tmp_17_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_9_b <= MUX1HOT_v_32_5_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_2_i_s_din_mxwt,
      twiddle_h_rsc_0_4_i_s_din_mxwt, twiddle_h_rsc_0_6_i_s_din_mxwt, twiddle_h_rsc_0_8_i_s_din_mxwt,
      STD_LOGIC_VECTOR'( (or_dcpl_29 OR INNER_LOOP1_tw_h_and_40_cse) & INNER_LOOP1_tw_h_and_41_cse
      & INNER_LOOP1_tw_h_and_42_cse & INNER_LOOP1_tw_h_and_43_cse & (fsm_output(8))));
  mult_t_mul_cmp_9_z <= mult_t_mul_cmp_9_z_1;

  mult_t_mul_cmp_10 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_10_a,
      b => mult_t_mul_cmp_10_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_10_z_1
    );
  mult_t_mul_cmp_10_a <= MUX1HOT_v_32_4_2(mult_t_mul_cmp_10_a_mx0w0, mult_t_mul_cmp_10_a_mx0w3,
      mult_t_mul_cmp_10_a_mx0w2, tmp_19_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_10_b <= MUX1HOT_v_32_6_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_1_i_s_din_mxwt,
      twiddle_h_rsc_0_4_i_s_din_mxwt, twiddle_h_rsc_0_5_i_s_din_mxwt, twiddle_h_rsc_0_9_i_s_din_mxwt,
      twiddle_h_rsc_0_8_i_s_din_mxwt, STD_LOGIC_VECTOR'( INNER_LOOP1_tw_h_or_1_cse
      & INNER_LOOP1_tw_h_and_37_cse & INNER_LOOP1_tw_h_and_38_cse & INNER_LOOP1_tw_h_and_39_cse
      & or_tmp_806 & and_1929_cse));
  mult_t_mul_cmp_10_z <= mult_t_mul_cmp_10_z_1;

  mult_t_mul_cmp_11 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_11_a,
      b => mult_t_mul_cmp_11_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_11_z_1
    );
  mult_t_mul_cmp_11_a <= MUX1HOT_v_32_4_2(mult_t_mul_cmp_11_a_mx0w0, mult_t_mul_cmp_11_a_mx0w3,
      mult_t_mul_cmp_11_a_mx0w2, tmp_21_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_11_b <= MUX1HOT_v_32_4_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_4_i_s_din_mxwt,
      twiddle_h_rsc_0_10_i_s_din_mxwt, twiddle_h_rsc_0_8_i_s_din_mxwt, STD_LOGIC_VECTOR'(
      (and_1948_cse OR or_dcpl_29) & or_tmp_812 & or_tmp_814 & and_1944_cse));
  mult_t_mul_cmp_11_z <= mult_t_mul_cmp_11_z_1;

  mult_t_mul_cmp_12 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_12_a,
      b => mult_t_mul_cmp_12_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_12_z_1
    );
  mult_t_mul_cmp_12_a <= mult_4_t_mux1h_rmff;
  mult_t_mul_cmp_12_b <= MUX1HOT_v_32_8_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_1_i_s_din_mxwt,
      twiddle_h_rsc_0_2_i_s_din_mxwt, twiddle_h_rsc_0_3_i_s_din_mxwt, twiddle_h_rsc_0_8_i_s_din_mxwt,
      twiddle_h_rsc_0_9_i_s_din_mxwt, twiddle_h_rsc_0_10_i_s_din_mxwt, twiddle_h_rsc_0_11_i_s_din_mxwt,
      STD_LOGIC_VECTOR'( INNER_LOOP1_tw_h_or_cse & INNER_LOOP1_tw_h_and_30_cse &
      INNER_LOOP1_tw_h_and_31_cse & INNER_LOOP1_tw_h_and_32_cse & INNER_LOOP1_tw_h_and_49_cse
      & INNER_LOOP1_tw_h_and_51_cse & INNER_LOOP1_tw_h_and_53_cse & INNER_LOOP1_tw_h_and_55_cse));
  mult_t_mul_cmp_12_z <= mult_t_mul_cmp_12_z_1;

  mult_t_mul_cmp_13 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_13_a,
      b => mult_t_mul_cmp_13_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_13_z_1
    );
  mult_t_mul_cmp_13_a <= MUX1HOT_v_32_4_2(mult_t_mul_cmp_13_a_mx0w0, tmp_7_lpi_3_dfm_mx0,
      mult_t_mul_cmp_13_a_mx0w2, tmp_25_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_13_b <= MUX1HOT_v_32_3_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_2_i_s_din_mxwt,
      twiddle_h_rsc_0_12_i_s_din_mxwt, STD_LOGIC_VECTOR'( or_tmp_888 & or_tmp_827
      & (fsm_output(8))));
  mult_t_mul_cmp_13_z <= mult_t_mul_cmp_13_z_1;

  mult_t_mul_cmp_14 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_14_a,
      b => mult_t_mul_cmp_14_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_14_z_1
    );
  mult_t_mul_cmp_14_a <= MUX1HOT_v_32_4_2(mult_t_mul_cmp_14_a_mx0w0, tmp_5_lpi_3_dfm_mx0,
      mult_t_mul_cmp_14_a_mx0w2, tmp_27_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_14_b <= MUX1HOT_v_32_4_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_1_i_s_din_mxwt,
      twiddle_h_rsc_0_13_i_s_din_mxwt, twiddle_h_rsc_0_12_i_s_din_mxwt, STD_LOGIC_VECTOR'(
      or_tmp_895 & or_tmp_835 & or_tmp_806 & and_1929_cse));
  mult_t_mul_cmp_14_z <= mult_t_mul_cmp_14_z_1;

  mult_t_mul_cmp_15 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 52,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_t_mul_cmp_15_a,
      b => mult_t_mul_cmp_15_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_t_mul_cmp_15_z_1
    );
  mult_t_mul_cmp_15_a <= MUX1HOT_v_32_4_2(mult_t_mul_cmp_15_a_mx0w0, tmp_3_lpi_3_dfm_mx0,
      mult_t_mul_cmp_15_a_mx0w2, tmp_29_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_t_mul_cmp_15_b <= MUX1HOT_v_32_3_2(twiddle_h_rsc_0_0_i_s_din_mxwt, twiddle_h_rsc_0_14_i_s_din_mxwt,
      twiddle_h_rsc_0_12_i_s_din_mxwt, STD_LOGIC_VECTOR'( (or_dcpl_29 OR (fsm_output(6)))
      & or_tmp_814 & and_1944_cse));
  mult_t_mul_cmp_15_z <= mult_t_mul_cmp_15_z_1;

  mult_z_mul_cmp : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_a,
      b => mult_z_mul_cmp_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_z_1
    );
  mult_z_mul_cmp_a <= MUX1HOT_v_32_3_2(tmp_65_lpi_3_dfm_mx0, tmp_1_lpi_3_dfm_mx0,
      mult_t_mul_cmp_a_mx0w2, STD_LOGIC_VECTOR'( (fsm_output(2)) & c_or_cse & (fsm_output(6))));
  mult_z_mul_cmp_b <= MUX1HOT_v_32_9_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_8_i_s_din_mxwt,
      twiddle_rsc_0_9_i_s_din_mxwt, twiddle_rsc_0_10_i_s_din_mxwt, twiddle_rsc_0_11_i_s_din_mxwt,
      twiddle_rsc_0_12_i_s_din_mxwt, twiddle_rsc_0_13_i_s_din_mxwt, twiddle_rsc_0_14_i_s_din_mxwt,
      twiddle_rsc_0_15_i_s_din_mxwt, STD_LOGIC_VECTOR'( (NOT (fsm_output(6))) & INNER_LOOP1_tw_h_and_44_cse
      & INNER_LOOP1_tw_h_and_45_cse & INNER_LOOP1_tw_h_and_46_cse & INNER_LOOP1_tw_h_and_47_cse
      & INNER_LOOP1_tw_h_and_48_cse & INNER_LOOP1_tw_h_and_50_cse & INNER_LOOP1_tw_h_and_52_cse
      & INNER_LOOP1_tw_h_and_54_cse));
  mult_z_mul_cmp_z <= mult_z_mul_cmp_z_1;

  mult_z_mul_cmp_1 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_1_a,
      b => mult_z_mul_cmp_1_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_1_z_1
    );
  mult_z_mul_cmp_1_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_1_z(51 DOWNTO 20)), (mult_t_mul_cmp_11_z(51
      DOWNTO 20)), (mult_t_mul_cmp_12_z(51 DOWNTO 20)), STD_LOGIC_VECTOR'( or_dcpl_29
      & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_1_b <= p_sva;
  mult_z_mul_cmp_1_z <= mult_z_mul_cmp_1_z_1;

  mult_z_mul_cmp_2 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_2_a,
      b => mult_z_mul_cmp_2_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_2_z_1
    );
  mult_z_mul_cmp_2_a <= MUX1HOT_v_32_4_2(mult_t_mul_cmp_1_a_mx0w0, tmp_31_lpi_3_dfm_mx0,
      mult_t_mul_cmp_15_a_mx0w2, tmp_17_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_2_b <= MUX_v_32_2_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_8_i_s_din_mxwt,
      fsm_output(8));
  mult_z_mul_cmp_2_z <= mult_z_mul_cmp_2_z_1;

  mult_z_mul_cmp_3 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_3_a,
      b => mult_z_mul_cmp_3_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_3_z_1
    );
  mult_z_mul_cmp_3_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_2_z(51 DOWNTO 20)), (mult_t_mul_cmp_5_z(51
      DOWNTO 20)), (mult_t_mul_cmp_6_z(51 DOWNTO 20)), STD_LOGIC_VECTOR'( or_dcpl_29
      & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_3_b <= p_sva;
  mult_z_mul_cmp_3_z <= mult_z_mul_cmp_3_z_1;

  mult_z_mul_cmp_4 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_4_a,
      b => mult_z_mul_cmp_4_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_4_z_1
    );
  mult_z_mul_cmp_4_a <= MUX1HOT_v_32_4_2(tmp_93_lpi_3_dfm_mx0, tmp_29_lpi_3_dfm_mx0,
      tmp_125_lpi_3_dfm_mx0, mult_t_mul_cmp_12_a_mx0w3, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_4_b <= MUX1HOT_v_32_6_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_8_i_s_din_mxwt,
      twiddle_rsc_0_10_i_s_din_mxwt, twiddle_rsc_0_12_i_s_din_mxwt, twiddle_rsc_0_14_i_s_din_mxwt,
      twiddle_rsc_0_4_i_s_din_mxwt, STD_LOGIC_VECTOR'( or_dcpl_29 & INNER_LOOP1_tw_h_and_40_cse
      & INNER_LOOP1_tw_h_and_41_cse & INNER_LOOP1_tw_h_and_42_cse & INNER_LOOP1_tw_h_and_43_cse
      & (fsm_output(8))));
  mult_z_mul_cmp_4_z <= mult_z_mul_cmp_4_z_1;

  mult_z_mul_cmp_5 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_5_a,
      b => mult_z_mul_cmp_5_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_5_z_1
    );
  mult_z_mul_cmp_5_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_3_z(51 DOWNTO 20)), (mult_t_mul_cmp_12_z(51
      DOWNTO 20)), (mult_t_mul_cmp_13_z(51 DOWNTO 20)), STD_LOGIC_VECTOR'( or_dcpl_29
      & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_5_b <= p_sva;
  mult_z_mul_cmp_5_z <= mult_z_mul_cmp_5_z_1;

  mult_z_mul_cmp_6 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_6_a,
      b => mult_z_mul_cmp_6_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_6_z_1
    );
  mult_z_mul_cmp_6_a <= MUX1HOT_v_32_4_2(tmp_91_lpi_3_dfm_mx0, tmp_27_lpi_3_dfm_mx0,
      mult_t_mul_cmp_8_a_mx0w2, tmp_31_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_6_b <= MUX1HOT_v_32_12_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_1_i_s_din_mxwt,
      twiddle_rsc_0_2_i_s_din_mxwt, twiddle_rsc_0_3_i_s_din_mxwt, twiddle_rsc_0_4_i_s_din_mxwt,
      twiddle_rsc_0_5_i_s_din_mxwt, twiddle_rsc_0_6_i_s_din_mxwt, twiddle_rsc_0_7_i_s_din_mxwt,
      twiddle_rsc_0_12_i_s_din_mxwt, twiddle_rsc_0_13_i_s_din_mxwt, twiddle_rsc_0_14_i_s_din_mxwt,
      twiddle_rsc_0_15_i_s_din_mxwt, STD_LOGIC_VECTOR'( INNER_LOOP1_tw_h_or_3_cse
      & INNER_LOOP1_tw_h_and_45_cse & INNER_LOOP1_tw_h_and_46_cse & INNER_LOOP1_tw_h_and_47_cse
      & INNER_LOOP1_tw_h_and_48_cse & INNER_LOOP1_tw_h_and_50_cse & INNER_LOOP1_tw_h_and_52_cse
      & INNER_LOOP1_tw_h_and_54_cse & INNER_LOOP1_tw_h_and_49_cse & INNER_LOOP1_tw_h_and_51_cse
      & INNER_LOOP1_tw_h_and_53_cse & INNER_LOOP1_tw_h_and_55_cse));
  mult_z_mul_cmp_6_z <= mult_z_mul_cmp_6_z_1;

  mult_z_mul_cmp_7 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_7_a,
      b => mult_z_mul_cmp_7_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_7_z_1
    );
  mult_z_mul_cmp_7_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_4_z(51 DOWNTO 20)), (mult_t_mul_cmp_2_z(51
      DOWNTO 20)), (mult_t_mul_cmp_3_z(51 DOWNTO 20)), STD_LOGIC_VECTOR'( or_dcpl_29
      & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_7_b <= p_sva;
  mult_z_mul_cmp_7_z <= mult_z_mul_cmp_7_z_1;

  mult_z_mul_cmp_8 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_8_a,
      b => mult_z_mul_cmp_8_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_8_z_1
    );
  mult_z_mul_cmp_8_a <= MUX1HOT_v_32_4_2(tmp_89_lpi_3_dfm_mx0, tmp_25_lpi_3_dfm_mx0,
      mult_t_mul_cmp_14_a_mx0w2, tmp_19_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_8_b <= MUX1HOT_v_32_4_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_1_i_s_din_mxwt,
      twiddle_rsc_0_9_i_s_din_mxwt, twiddle_rsc_0_8_i_s_din_mxwt, STD_LOGIC_VECTOR'(
      or_tmp_895 & or_tmp_835 & or_tmp_806 & and_1929_cse));
  mult_z_mul_cmp_8_z <= mult_z_mul_cmp_8_z_1;

  mult_z_mul_cmp_9 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_9_a,
      b => mult_z_mul_cmp_9_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_9_z_1
    );
  mult_z_mul_cmp_9_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_5_z(51 DOWNTO 20)), (mult_t_mul_cmp_10_z(51
      DOWNTO 20)), (mult_t_mul_cmp_11_z(51 DOWNTO 20)), STD_LOGIC_VECTOR'( or_dcpl_29
      & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_9_b <= p_sva;
  mult_z_mul_cmp_9_z <= mult_z_mul_cmp_9_z_1;

  mult_z_mul_cmp_10 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_10_a,
      b => mult_z_mul_cmp_10_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_10_z_1
    );
  mult_z_mul_cmp_10_a <= MUX1HOT_v_32_4_2(tmp_87_lpi_3_dfm_mx0, tmp_23_lpi_3_dfm_mx0,
      mult_t_mul_cmp_7_a_mx0w2, mult_t_mul_cmp_9_a_mx0w3, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_10_b <= MUX1HOT_v_32_6_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_8_i_s_din_mxwt,
      twiddle_rsc_0_4_i_s_din_mxwt, twiddle_rsc_0_5_i_s_din_mxwt, twiddle_rsc_0_6_i_s_din_mxwt,
      twiddle_rsc_0_7_i_s_din_mxwt, STD_LOGIC_VECTOR'( or_dcpl_29 & (fsm_output(6))
      & INNER_LOOP1_tw_h_and_49_cse & INNER_LOOP1_tw_h_and_51_cse & INNER_LOOP1_tw_h_and_53_cse
      & INNER_LOOP1_tw_h_and_55_cse));
  mult_z_mul_cmp_10_z <= mult_z_mul_cmp_10_z_1;

  mult_z_mul_cmp_11 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_11_a,
      b => mult_z_mul_cmp_11_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_11_z_1
    );
  mult_z_mul_cmp_11_a <= MUX_v_32_2_2((mult_t_mul_cmp_6_z(51 DOWNTO 20)), (mult_t_mul_cmp_7_z(51
      DOWNTO 20)), fsm_output(8));
  mult_z_mul_cmp_11_b <= p_sva;
  mult_z_mul_cmp_11_z <= mult_z_mul_cmp_11_z_1;

  mult_z_mul_cmp_12 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_12_a,
      b => mult_z_mul_cmp_12_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_12_z_1
    );
  mult_z_mul_cmp_12_a <= MUX1HOT_v_32_4_2(tmp_85_lpi_3_dfm_mx0, tmp_21_lpi_3_dfm_mx0,
      mult_t_mul_cmp_13_a_mx0w2, tmp_7_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_12_b <= MUX1HOT_v_32_4_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_2_i_s_din_mxwt,
      twiddle_rsc_0_1_i_s_din_mxwt, twiddle_rsc_0_3_i_s_din_mxwt, STD_LOGIC_VECTOR'(
      (or_tmp_888 OR INNER_LOOP1_tw_h_and_49_cse) & (or_tmp_827 OR INNER_LOOP1_tw_h_and_53_cse)
      & INNER_LOOP1_tw_h_and_51_cse & INNER_LOOP1_tw_h_and_55_cse));
  mult_z_mul_cmp_12_z <= mult_z_mul_cmp_12_z_1;

  mult_z_mul_cmp_13 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_13_a,
      b => mult_z_mul_cmp_13_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_13_z_1
    );
  mult_z_mul_cmp_13_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_7_z(51 DOWNTO 20)), (mult_t_mul_cmp_1_z(51
      DOWNTO 20)), (mult_t_mul_cmp_2_z(51 DOWNTO 20)), STD_LOGIC_VECTOR'( or_dcpl_29
      & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_13_b <= p_sva;
  mult_z_mul_cmp_13_z <= mult_z_mul_cmp_13_z_1;

  mult_z_mul_cmp_14 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_14_a,
      b => mult_z_mul_cmp_14_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_14_z_1
    );
  mult_z_mul_cmp_14_a <= MUX1HOT_v_32_4_2(tmp_83_lpi_3_dfm_mx0, tmp_19_lpi_3_dfm_mx0,
      mult_t_mul_cmp_2_a_mx0w2, tmp_29_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_14_b <= MUX1HOT_v_32_6_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_8_i_s_din_mxwt,
      twiddle_rsc_0_9_i_s_din_mxwt, twiddle_rsc_0_12_i_s_din_mxwt, twiddle_rsc_0_13_i_s_din_mxwt,
      twiddle_rsc_0_14_i_s_din_mxwt, STD_LOGIC_VECTOR'( or_dcpl_29 & INNER_LOOP1_tw_h_and_36_cse
      & INNER_LOOP1_tw_h_and_37_cse & (INNER_LOOP1_tw_h_and_38_cse OR and_1944_cse)
      & INNER_LOOP1_tw_h_and_39_cse & or_tmp_814));
  mult_z_mul_cmp_14_z <= mult_z_mul_cmp_14_z_1;

  mult_z_mul_cmp_15 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_15_a,
      b => mult_z_mul_cmp_15_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_15_z_1
    );
  mult_z_mul_cmp_15_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_8_z(51 DOWNTO 20)), (mult_t_mul_cmp_13_z(51
      DOWNTO 20)), (mult_t_mul_cmp_14_z(51 DOWNTO 20)), STD_LOGIC_VECTOR'( or_dcpl_29
      & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_15_b <= p_sva;
  mult_z_mul_cmp_15_z <= mult_z_mul_cmp_15_z_1;

  mult_z_mul_cmp_16 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_16_a,
      b => mult_z_mul_cmp_16_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_16_z_1
    );
  mult_z_mul_cmp_16_a <= MUX1HOT_v_32_4_2(tmp_81_lpi_3_dfm_mx0, tmp_17_lpi_3_dfm_mx0,
      mult_t_mul_cmp_9_a_mx0w2, tmp_3_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_16_b <= MUX1HOT_v_32_5_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_2_i_s_din_mxwt,
      twiddle_rsc_0_4_i_s_din_mxwt, twiddle_rsc_0_6_i_s_din_mxwt, twiddle_rsc_0_1_i_s_din_mxwt,
      STD_LOGIC_VECTOR'( (or_tmp_804 OR INNER_LOOP1_tw_h_and_40_cse) & INNER_LOOP1_tw_h_and_41_cse
      & INNER_LOOP1_tw_h_and_42_cse & INNER_LOOP1_tw_h_and_43_cse & or_tmp_806));
  mult_z_mul_cmp_16_z <= mult_z_mul_cmp_16_z_1;

  mult_z_mul_cmp_17 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_17_a,
      b => mult_z_mul_cmp_17_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_17_z_1
    );
  mult_z_mul_cmp_17_a <= MUX_v_32_2_2((mult_t_mul_cmp_9_z(51 DOWNTO 20)), (mult_t_mul_cmp_10_z(51
      DOWNTO 20)), fsm_output(8));
  mult_z_mul_cmp_17_b <= p_sva;
  mult_z_mul_cmp_17_z <= mult_z_mul_cmp_17_z_1;

  mult_z_mul_cmp_18 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_18_a,
      b => mult_z_mul_cmp_18_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_18_z_1
    );
  mult_z_mul_cmp_18_a <= MUX1HOT_v_32_4_2(mult_t_mul_cmp_9_a_mx0w0, mult_t_mul_cmp_9_a_mx0w3,
      mult_t_mul_cmp_6_a_mx0w2, tmp_21_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_18_b <= MUX1HOT_v_32_4_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_9_i_s_din_mxwt,
      twiddle_rsc_0_8_i_s_din_mxwt, twiddle_rsc_0_10_i_s_din_mxwt, STD_LOGIC_VECTOR'(
      or_dcpl_29 & or_tmp_835 & (and_1994_cse OR and_1944_cse) & or_tmp_814));
  mult_z_mul_cmp_18_z <= mult_z_mul_cmp_18_z_1;

  mult_z_mul_cmp_19 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_19_a,
      b => mult_z_mul_cmp_19_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_19_z_1
    );
  mult_z_mul_cmp_19_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_10_z(51 DOWNTO 20)), (mult_t_mul_cmp_4_z(51
      DOWNTO 20)), (mult_t_mul_cmp_5_z(51 DOWNTO 20)), STD_LOGIC_VECTOR'( or_dcpl_29
      & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_19_b <= p_sva;
  mult_z_mul_cmp_19_z <= mult_z_mul_cmp_19_z_1;

  mult_z_mul_cmp_20 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_20_a,
      b => mult_z_mul_cmp_20_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_20_z_1
    );
  mult_z_mul_cmp_20_a <= MUX1HOT_v_32_4_2(mult_t_mul_cmp_10_a_mx0w0, mult_t_mul_cmp_10_a_mx0w3,
      tmp_121_lpi_3_dfm_mx0, mult_t_mul_cmp_11_a_mx0w3, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_20_b <= MUX1HOT_v_32_5_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_12_i_s_din_mxwt,
      twiddle_rsc_0_8_i_s_din_mxwt, twiddle_rsc_0_5_i_s_din_mxwt, twiddle_rsc_0_4_i_s_din_mxwt,
      STD_LOGIC_VECTOR'( or_dcpl_29 & or_tmp_812 & and_1948_cse & or_tmp_806 & and_1929_cse));
  mult_z_mul_cmp_20_z <= mult_z_mul_cmp_20_z_1;

  mult_z_mul_cmp_21 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_21_a,
      b => mult_z_mul_cmp_21_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_21_z_1
    );
  mult_z_mul_cmp_21_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_11_z(51 DOWNTO 20)), (mult_t_mul_cmp_14_z(51
      DOWNTO 20)), (mult_t_mul_cmp_15_z(51 DOWNTO 20)), STD_LOGIC_VECTOR'( or_dcpl_29
      & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_21_b <= p_sva;
  mult_z_mul_cmp_21_z <= mult_z_mul_cmp_21_z_1;

  mult_z_mul_cmp_22 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_22_a,
      b => mult_z_mul_cmp_22_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_22_z_1
    );
  mult_z_mul_cmp_22_a <= MUX1HOT_v_32_4_2(mult_t_mul_cmp_11_a_mx0w0, mult_t_mul_cmp_11_a_mx0w3,
      mult_t_mul_cmp_10_a_mx0w2, tmp_27_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_22_b <= MUX1HOT_v_32_6_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_1_i_s_din_mxwt,
      twiddle_rsc_0_4_i_s_din_mxwt, twiddle_rsc_0_5_i_s_din_mxwt, twiddle_rsc_0_13_i_s_din_mxwt,
      twiddle_rsc_0_12_i_s_din_mxwt, STD_LOGIC_VECTOR'( INNER_LOOP1_tw_h_or_1_cse
      & INNER_LOOP1_tw_h_and_37_cse & INNER_LOOP1_tw_h_and_38_cse & INNER_LOOP1_tw_h_and_39_cse
      & or_tmp_806 & and_1929_cse));
  mult_z_mul_cmp_22_z <= mult_z_mul_cmp_22_z_1;

  mult_z_mul_cmp_23 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_23_a,
      b => mult_z_mul_cmp_23_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_23_z_1
    );
  mult_z_mul_cmp_23_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_12_z(51 DOWNTO 20)), (mult_t_mul_cmp_3_z(51
      DOWNTO 20)), (mult_t_mul_cmp_4_z(51 DOWNTO 20)), STD_LOGIC_VECTOR'( or_dcpl_29
      & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_23_b <= p_sva;
  mult_z_mul_cmp_23_z <= mult_z_mul_cmp_23_z_1;

  mult_z_mul_cmp_24 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_24_a,
      b => mult_z_mul_cmp_24_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_24_z_1
    );
  mult_z_mul_cmp_24_a <= mult_4_t_mux1h_rmff;
  mult_z_mul_cmp_24_b <= MUX1HOT_v_32_8_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_1_i_s_din_mxwt,
      twiddle_rsc_0_2_i_s_din_mxwt, twiddle_rsc_0_3_i_s_din_mxwt, twiddle_rsc_0_8_i_s_din_mxwt,
      twiddle_rsc_0_9_i_s_din_mxwt, twiddle_rsc_0_10_i_s_din_mxwt, twiddle_rsc_0_11_i_s_din_mxwt,
      STD_LOGIC_VECTOR'( INNER_LOOP1_tw_h_or_cse & INNER_LOOP1_tw_h_and_30_cse &
      INNER_LOOP1_tw_h_and_31_cse & INNER_LOOP1_tw_h_and_32_cse & INNER_LOOP1_tw_h_and_49_cse
      & INNER_LOOP1_tw_h_and_51_cse & INNER_LOOP1_tw_h_and_53_cse & INNER_LOOP1_tw_h_and_55_cse));
  mult_z_mul_cmp_24_z <= mult_z_mul_cmp_24_z_1;

  mult_z_mul_cmp_25 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_25_a,
      b => mult_z_mul_cmp_25_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_25_z_1
    );
  mult_z_mul_cmp_25_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_13_z(51 DOWNTO 20)), (mult_t_mul_cmp_8_z(51
      DOWNTO 20)), (mult_t_mul_cmp_9_z(51 DOWNTO 20)), STD_LOGIC_VECTOR'( or_dcpl_29
      & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_25_b <= p_sva;
  mult_z_mul_cmp_25_z <= mult_z_mul_cmp_25_z_1;

  mult_z_mul_cmp_26 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_26_a,
      b => mult_z_mul_cmp_26_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_26_z_1
    );
  mult_z_mul_cmp_26_a <= MUX1HOT_v_32_4_2(mult_t_mul_cmp_13_a_mx0w0, tmp_7_lpi_3_dfm_mx0,
      mult_t_mul_cmp_5_a_mx0w2, mult_t_mul_cmp_10_a_mx0w3, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_26_b <= MUX1HOT_v_32_5_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_10_i_s_din_mxwt,
      twiddle_rsc_0_8_i_s_din_mxwt, twiddle_rsc_0_6_i_s_din_mxwt, twiddle_rsc_0_4_i_s_din_mxwt,
      STD_LOGIC_VECTOR'( or_dcpl_29 & or_tmp_827 & and_1978_cse & or_tmp_814 & and_1944_cse));
  mult_z_mul_cmp_26_z <= mult_z_mul_cmp_26_z_1;

  mult_z_mul_cmp_27 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_27_a,
      b => mult_z_mul_cmp_27_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_27_z_1
    );
  mult_z_mul_cmp_27_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_14_z(51 DOWNTO 20)), (mult_t_mul_cmp_7_z(51
      DOWNTO 20)), (mult_t_mul_cmp_8_z(51 DOWNTO 20)), STD_LOGIC_VECTOR'( or_dcpl_29
      & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_27_b <= p_sva;
  mult_z_mul_cmp_27_z <= mult_z_mul_cmp_27_z_1;

  mult_z_mul_cmp_28 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_28_a,
      b => mult_z_mul_cmp_28_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_28_z_1
    );
  mult_z_mul_cmp_28_a <= MUX1HOT_v_32_3_2(mult_t_mul_cmp_14_a_mx0w0, tmp_5_lpi_3_dfm_mx0,
      mult_t_mul_cmp_11_a_mx0w2, STD_LOGIC_VECTOR'( (fsm_output(2)) & c_or_cse &
      (fsm_output(6))));
  mult_z_mul_cmp_28_b <= MUX1HOT_v_32_3_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_4_i_s_din_mxwt,
      twiddle_rsc_0_2_i_s_din_mxwt, STD_LOGIC_VECTOR'( (and_1948_cse OR or_dcpl_29
      OR and_1944_cse) & or_tmp_812 & or_tmp_814));
  mult_z_mul_cmp_28_z <= mult_z_mul_cmp_28_z_1;

  mult_z_mul_cmp_29 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_29_a,
      b => mult_z_mul_cmp_29_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_29_z_1
    );
  mult_z_mul_cmp_29_a <= MUX1HOT_v_32_3_2((mult_t_mul_cmp_15_z(51 DOWNTO 20)), (mult_t_mul_cmp_z(51
      DOWNTO 20)), (mult_t_mul_cmp_1_z(51 DOWNTO 20)), STD_LOGIC_VECTOR'( or_dcpl_29
      & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_29_b <= p_sva;
  mult_z_mul_cmp_29_z <= mult_z_mul_cmp_29_z_1;

  mult_z_mul_cmp_30 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_30_a,
      b => mult_z_mul_cmp_30_b,
      clk => clk,
      en => mult_t_mul_cmp_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_30_z_1
    );
  mult_z_mul_cmp_30_a <= MUX1HOT_v_32_4_2(mult_t_mul_cmp_15_a_mx0w0, tmp_3_lpi_3_dfm_mx0,
      mult_t_mul_cmp_4_a_mx0w2, tmp_25_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  mult_z_mul_cmp_30_b <= MUX1HOT_v_32_6_2(twiddle_rsc_0_0_i_s_din_mxwt, twiddle_rsc_0_8_i_s_din_mxwt,
      twiddle_rsc_0_9_i_s_din_mxwt, twiddle_rsc_0_10_i_s_din_mxwt, twiddle_rsc_0_11_i_s_din_mxwt,
      twiddle_rsc_0_12_i_s_din_mxwt, STD_LOGIC_VECTOR'( or_dcpl_29 & INNER_LOOP1_tw_h_and_29_cse
      & INNER_LOOP1_tw_h_and_30_cse & INNER_LOOP1_tw_h_and_31_cse & INNER_LOOP1_tw_h_and_32_cse
      & (fsm_output(8))));
  mult_z_mul_cmp_30_z <= mult_z_mul_cmp_30_z_1;

  mult_z_mul_cmp_31 : work.mgc_comps.mgc_mul_pipe
    GENERIC MAP(
      width_a => 32,
      signd_a => 0,
      width_b => 32,
      signd_b => 0,
      width_z => 32,
      clock_edge => 1,
      enable_active => 1,
      a_rst_active => 0,
      s_rst_active => 1,
      stages => 2,
      n_inreg => 2
      )
    PORT MAP(
      a => mult_z_mul_cmp_31_a,
      b => mult_z_mul_cmp_31_b,
      clk => clk,
      en => mult_z_mul_cmp_1_en,
      a_rst => '1',
      s_rst => rst,
      z => mult_z_mul_cmp_31_z_1
    );
  mult_z_mul_cmp_31_a <= MUX_v_32_2_2((mult_t_mul_cmp_z(51 DOWNTO 20)), (mult_t_mul_cmp_15_z(51
      DOWNTO 20)), fsm_output(6));
  mult_z_mul_cmp_31_b <= p_sva;
  mult_z_mul_cmp_31_z <= mult_z_mul_cmp_31_z_1;

  operator_33_true_3_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_bl_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 1,
      width_s => 3,
      width_z => 2
      )
    PORT MAP(
      a => operator_33_true_3_lshift_rg_a,
      s => operator_33_true_3_lshift_rg_s,
      z => operator_33_true_3_lshift_rg_z
    );
  operator_33_true_3_lshift_rg_a(0) <= '1';
  operator_33_true_3_lshift_rg_s <= STD_LOGIC_VECTOR'( '0' & (NOT c_1_sva_1) & '0');
  operator_33_true_3_lshift_psp_1_0_sva_mx0w2 <= operator_33_true_3_lshift_rg_z;

  operator_33_true_1_lshift_rg : work.mgc_shift_comps_v5.mgc_shift_l_v5
    GENERIC MAP(
      width_a => 1,
      signd_a => 1,
      width_s => 4,
      width_z => 9
      )
    PORT MAP(
      a => operator_33_true_1_lshift_rg_a,
      s => operator_33_true_1_lshift_rg_s,
      z => operator_33_true_1_lshift_rg_z
    );
  operator_33_true_1_lshift_rg_a(0) <= '1';
  operator_33_true_1_lshift_rg_s <= (MUX1HOT_v_3_3_2(operator_20_false_acc_cse_sva_mx0w0,
      operator_20_false_acc_cse_sva, (STD_LOGIC_VECTOR'( "00") & (NOT c_1_sva_1)),
      STD_LOGIC_VECTOR'( (fsm_output(1)) & (fsm_output(3)) & (fsm_output(5))))) &
      ((NOT (fsm_output(3))) OR (fsm_output(1)) OR (fsm_output(5)));
  z_out_32 <= operator_33_true_1_lshift_rg_z;

  peaseNTT_core_wait_dp_inst : peaseNTT_core_wait_dp
    PORT MAP(
      yt_rsc_0_0_cgo_iro => or_67_rmff,
      yt_rsc_0_0_i_clken_d => yt_rsc_0_0_i_clken_d,
      yt_rsc_0_16_cgo_iro => or_166_rmff,
      yt_rsc_0_16_i_clken_d => yt_rsc_0_16_i_clken_d,
      yt_rsc_1_0_cgo_iro => or_248_rmff,
      yt_rsc_1_0_i_clken_d => yt_rsc_1_0_i_clken_d,
      yt_rsc_1_16_cgo_iro => or_347_rmff,
      yt_rsc_1_16_i_clken_d => yt_rsc_1_16_i_clken_d,
      ensig_cgo_iro => or_833_rmff,
      ensig_cgo_iro_17 => or_956_rmff,
      core_wen => core_wen,
      yt_rsc_0_0_cgo => reg_yt_rsc_0_0_cgo_cse,
      yt_rsc_0_16_cgo => reg_yt_rsc_0_16_cgo_cse,
      yt_rsc_1_0_cgo => reg_yt_rsc_1_0_cgo_cse,
      yt_rsc_1_16_cgo => reg_yt_rsc_1_16_cgo_cse,
      ensig_cgo => reg_ensig_cgo_cse,
      mult_t_mul_cmp_en => mult_t_mul_cmp_en,
      ensig_cgo_17 => reg_ensig_cgo_17_cse,
      mult_z_mul_cmp_1_en => mult_z_mul_cmp_1_en
    );
  peaseNTT_core_xt_rsc_0_0_i_1_inst : peaseNTT_core_xt_rsc_0_0_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_0_i_qa_d => peaseNTT_core_xt_rsc_0_0_i_1_inst_xt_rsc_0_0_i_qa_d,
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      xt_rsc_0_0_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      core_wten => core_wten,
      xt_rsc_0_0_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_0_i_1_inst_xt_rsc_0_0_i_qa_d_mxwt,
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_0_i_wea_d_pff => xt_rsc_0_0_i_wea_d_iff,
      xt_rsc_0_0_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_0_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_0_i_1_inst_xt_rsc_0_0_i_qa_d <= xt_rsc_0_0_i_qa_d;
  xt_rsc_0_0_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_0_i_1_inst_xt_rsc_0_0_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_1_i_1_inst : peaseNTT_core_xt_rsc_0_1_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_1_i_qa_d => peaseNTT_core_xt_rsc_0_1_i_1_inst_xt_rsc_0_1_i_qa_d,
      xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_1_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_1_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_1_i_1_inst_xt_rsc_0_1_i_qa_d_mxwt,
      xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_1_i_wea_d_pff => xt_rsc_0_1_i_wea_d_iff,
      xt_rsc_0_1_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_1_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_1_i_1_inst_xt_rsc_0_1_i_qa_d <= xt_rsc_0_1_i_qa_d;
  xt_rsc_0_1_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_1_i_1_inst_xt_rsc_0_1_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_2_i_1_inst : peaseNTT_core_xt_rsc_0_2_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_2_i_qa_d => peaseNTT_core_xt_rsc_0_2_i_1_inst_xt_rsc_0_2_i_qa_d,
      xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_2_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_2_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_2_i_1_inst_xt_rsc_0_2_i_qa_d_mxwt,
      xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_2_i_wea_d_pff => xt_rsc_0_2_i_wea_d_iff,
      xt_rsc_0_2_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_2_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_2_i_1_inst_xt_rsc_0_2_i_qa_d <= xt_rsc_0_2_i_qa_d;
  xt_rsc_0_2_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_2_i_1_inst_xt_rsc_0_2_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_3_i_1_inst : peaseNTT_core_xt_rsc_0_3_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_3_i_qa_d => peaseNTT_core_xt_rsc_0_3_i_1_inst_xt_rsc_0_3_i_qa_d,
      xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_3_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_3_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_3_i_1_inst_xt_rsc_0_3_i_qa_d_mxwt,
      xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_3_i_wea_d_pff => xt_rsc_0_3_i_wea_d_iff,
      xt_rsc_0_3_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_3_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_3_i_1_inst_xt_rsc_0_3_i_qa_d <= xt_rsc_0_3_i_qa_d;
  xt_rsc_0_3_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_3_i_1_inst_xt_rsc_0_3_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_4_i_1_inst : peaseNTT_core_xt_rsc_0_4_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_4_i_qa_d => peaseNTT_core_xt_rsc_0_4_i_1_inst_xt_rsc_0_4_i_qa_d,
      xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_4_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_4_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_4_i_1_inst_xt_rsc_0_4_i_qa_d_mxwt,
      xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_4_i_wea_d_pff => xt_rsc_0_4_i_wea_d_iff,
      xt_rsc_0_4_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_4_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_4_i_1_inst_xt_rsc_0_4_i_qa_d <= xt_rsc_0_4_i_qa_d;
  xt_rsc_0_4_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_4_i_1_inst_xt_rsc_0_4_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_5_i_1_inst : peaseNTT_core_xt_rsc_0_5_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_5_i_qa_d => peaseNTT_core_xt_rsc_0_5_i_1_inst_xt_rsc_0_5_i_qa_d,
      xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_5_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_5_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_5_i_1_inst_xt_rsc_0_5_i_qa_d_mxwt,
      xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_5_i_wea_d_pff => xt_rsc_0_5_i_wea_d_iff,
      xt_rsc_0_5_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_5_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_5_i_1_inst_xt_rsc_0_5_i_qa_d <= xt_rsc_0_5_i_qa_d;
  xt_rsc_0_5_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_5_i_1_inst_xt_rsc_0_5_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_6_i_1_inst : peaseNTT_core_xt_rsc_0_6_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_6_i_qa_d => peaseNTT_core_xt_rsc_0_6_i_1_inst_xt_rsc_0_6_i_qa_d,
      xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_6_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_6_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_6_i_1_inst_xt_rsc_0_6_i_qa_d_mxwt,
      xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_6_i_wea_d_pff => xt_rsc_0_6_i_wea_d_iff,
      xt_rsc_0_6_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_6_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_6_i_1_inst_xt_rsc_0_6_i_qa_d <= xt_rsc_0_6_i_qa_d;
  xt_rsc_0_6_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_6_i_1_inst_xt_rsc_0_6_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_7_i_1_inst : peaseNTT_core_xt_rsc_0_7_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_7_i_qa_d => peaseNTT_core_xt_rsc_0_7_i_1_inst_xt_rsc_0_7_i_qa_d,
      xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_7_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_7_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_7_i_1_inst_xt_rsc_0_7_i_qa_d_mxwt,
      xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_7_i_wea_d_pff => xt_rsc_0_7_i_wea_d_iff,
      xt_rsc_0_7_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_7_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_7_i_1_inst_xt_rsc_0_7_i_qa_d <= xt_rsc_0_7_i_qa_d;
  xt_rsc_0_7_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_7_i_1_inst_xt_rsc_0_7_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_8_i_1_inst : peaseNTT_core_xt_rsc_0_8_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_8_i_qa_d => peaseNTT_core_xt_rsc_0_8_i_1_inst_xt_rsc_0_8_i_qa_d,
      xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_8_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_8_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_8_i_1_inst_xt_rsc_0_8_i_qa_d_mxwt,
      xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_8_i_wea_d_pff => xt_rsc_0_8_i_wea_d_iff,
      xt_rsc_0_8_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_8_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_8_i_1_inst_xt_rsc_0_8_i_qa_d <= xt_rsc_0_8_i_qa_d;
  xt_rsc_0_8_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_8_i_1_inst_xt_rsc_0_8_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_9_i_1_inst : peaseNTT_core_xt_rsc_0_9_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_9_i_qa_d => peaseNTT_core_xt_rsc_0_9_i_1_inst_xt_rsc_0_9_i_qa_d,
      xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_9_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_9_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_9_i_1_inst_xt_rsc_0_9_i_qa_d_mxwt,
      xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_9_i_wea_d_pff => xt_rsc_0_9_i_wea_d_iff,
      xt_rsc_0_9_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_9_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_9_i_1_inst_xt_rsc_0_9_i_qa_d <= xt_rsc_0_9_i_qa_d;
  xt_rsc_0_9_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_9_i_1_inst_xt_rsc_0_9_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_10_i_1_inst : peaseNTT_core_xt_rsc_0_10_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_10_i_qa_d => peaseNTT_core_xt_rsc_0_10_i_1_inst_xt_rsc_0_10_i_qa_d,
      xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_10_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_10_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_10_i_1_inst_xt_rsc_0_10_i_qa_d_mxwt,
      xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_10_i_wea_d_pff => xt_rsc_0_10_i_wea_d_iff,
      xt_rsc_0_10_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_10_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_10_i_1_inst_xt_rsc_0_10_i_qa_d <= xt_rsc_0_10_i_qa_d;
  xt_rsc_0_10_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_10_i_1_inst_xt_rsc_0_10_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_11_i_1_inst : peaseNTT_core_xt_rsc_0_11_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_11_i_qa_d => peaseNTT_core_xt_rsc_0_11_i_1_inst_xt_rsc_0_11_i_qa_d,
      xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_11_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_11_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_11_i_1_inst_xt_rsc_0_11_i_qa_d_mxwt,
      xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_11_i_wea_d_pff => xt_rsc_0_11_i_wea_d_iff,
      xt_rsc_0_11_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_11_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_11_i_1_inst_xt_rsc_0_11_i_qa_d <= xt_rsc_0_11_i_qa_d;
  xt_rsc_0_11_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_11_i_1_inst_xt_rsc_0_11_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_12_i_1_inst : peaseNTT_core_xt_rsc_0_12_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_12_i_qa_d => peaseNTT_core_xt_rsc_0_12_i_1_inst_xt_rsc_0_12_i_qa_d,
      xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_12_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_12_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_12_i_1_inst_xt_rsc_0_12_i_qa_d_mxwt,
      xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_12_i_wea_d_pff => xt_rsc_0_12_i_wea_d_iff,
      xt_rsc_0_12_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_12_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_12_i_1_inst_xt_rsc_0_12_i_qa_d <= xt_rsc_0_12_i_qa_d;
  xt_rsc_0_12_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_12_i_1_inst_xt_rsc_0_12_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_13_i_1_inst : peaseNTT_core_xt_rsc_0_13_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_13_i_qa_d => peaseNTT_core_xt_rsc_0_13_i_1_inst_xt_rsc_0_13_i_qa_d,
      xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_13_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_13_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_13_i_1_inst_xt_rsc_0_13_i_qa_d_mxwt,
      xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_13_i_wea_d_pff => xt_rsc_0_13_i_wea_d_iff,
      xt_rsc_0_13_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_13_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_13_i_1_inst_xt_rsc_0_13_i_qa_d <= xt_rsc_0_13_i_qa_d;
  xt_rsc_0_13_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_13_i_1_inst_xt_rsc_0_13_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_14_i_1_inst : peaseNTT_core_xt_rsc_0_14_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_14_i_qa_d => peaseNTT_core_xt_rsc_0_14_i_1_inst_xt_rsc_0_14_i_qa_d,
      xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_14_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_14_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_14_i_1_inst_xt_rsc_0_14_i_qa_d_mxwt,
      xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_14_i_wea_d_pff => xt_rsc_0_14_i_wea_d_iff,
      xt_rsc_0_14_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_14_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_14_i_1_inst_xt_rsc_0_14_i_qa_d <= xt_rsc_0_14_i_qa_d;
  xt_rsc_0_14_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_14_i_1_inst_xt_rsc_0_14_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_15_i_1_inst : peaseNTT_core_xt_rsc_0_15_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_15_i_qa_d => peaseNTT_core_xt_rsc_0_15_i_1_inst_xt_rsc_0_15_i_qa_d,
      xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_15_i_oswt => reg_xt_rsc_0_0_i_oswt_cse,
      xt_rsc_0_15_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_15_i_1_inst_xt_rsc_0_15_i_qa_d_mxwt,
      xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_15_i_wea_d_pff => xt_rsc_0_15_i_wea_d_iff,
      xt_rsc_0_15_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_0_15_i_oswt_pff => or_429_rmff
    );
  peaseNTT_core_xt_rsc_0_15_i_1_inst_xt_rsc_0_15_i_qa_d <= xt_rsc_0_15_i_qa_d;
  xt_rsc_0_15_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_15_i_1_inst_xt_rsc_0_15_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_16_i_1_inst : peaseNTT_core_xt_rsc_0_16_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_16_i_qa_d => peaseNTT_core_xt_rsc_0_16_i_1_inst_xt_rsc_0_16_i_qa_d,
      xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_16_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_16_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_16_i_1_inst_xt_rsc_0_16_i_qa_d_mxwt,
      xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_16_i_wea_d_pff => xt_rsc_0_16_i_wea_d_iff,
      xt_rsc_0_16_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_16_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_16_i_1_inst_xt_rsc_0_16_i_qa_d <= xt_rsc_0_16_i_qa_d;
  xt_rsc_0_16_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_16_i_1_inst_xt_rsc_0_16_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_17_i_1_inst : peaseNTT_core_xt_rsc_0_17_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_17_i_qa_d => peaseNTT_core_xt_rsc_0_17_i_1_inst_xt_rsc_0_17_i_qa_d,
      xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_17_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_17_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_17_i_1_inst_xt_rsc_0_17_i_qa_d_mxwt,
      xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_17_i_wea_d_pff => xt_rsc_0_17_i_wea_d_iff,
      xt_rsc_0_17_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_17_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_17_i_1_inst_xt_rsc_0_17_i_qa_d <= xt_rsc_0_17_i_qa_d;
  xt_rsc_0_17_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_17_i_1_inst_xt_rsc_0_17_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_18_i_1_inst : peaseNTT_core_xt_rsc_0_18_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_18_i_qa_d => peaseNTT_core_xt_rsc_0_18_i_1_inst_xt_rsc_0_18_i_qa_d,
      xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_18_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_18_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_18_i_1_inst_xt_rsc_0_18_i_qa_d_mxwt,
      xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_18_i_wea_d_pff => xt_rsc_0_18_i_wea_d_iff,
      xt_rsc_0_18_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_18_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_18_i_1_inst_xt_rsc_0_18_i_qa_d <= xt_rsc_0_18_i_qa_d;
  xt_rsc_0_18_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_18_i_1_inst_xt_rsc_0_18_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_19_i_1_inst : peaseNTT_core_xt_rsc_0_19_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_19_i_qa_d => peaseNTT_core_xt_rsc_0_19_i_1_inst_xt_rsc_0_19_i_qa_d,
      xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_19_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_19_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_19_i_1_inst_xt_rsc_0_19_i_qa_d_mxwt,
      xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_19_i_wea_d_pff => xt_rsc_0_19_i_wea_d_iff,
      xt_rsc_0_19_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_19_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_19_i_1_inst_xt_rsc_0_19_i_qa_d <= xt_rsc_0_19_i_qa_d;
  xt_rsc_0_19_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_19_i_1_inst_xt_rsc_0_19_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_20_i_1_inst : peaseNTT_core_xt_rsc_0_20_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_20_i_qa_d => peaseNTT_core_xt_rsc_0_20_i_1_inst_xt_rsc_0_20_i_qa_d,
      xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_20_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_20_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_20_i_1_inst_xt_rsc_0_20_i_qa_d_mxwt,
      xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_20_i_wea_d_pff => xt_rsc_0_20_i_wea_d_iff,
      xt_rsc_0_20_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_20_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_20_i_1_inst_xt_rsc_0_20_i_qa_d <= xt_rsc_0_20_i_qa_d;
  xt_rsc_0_20_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_20_i_1_inst_xt_rsc_0_20_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_21_i_1_inst : peaseNTT_core_xt_rsc_0_21_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_21_i_qa_d => peaseNTT_core_xt_rsc_0_21_i_1_inst_xt_rsc_0_21_i_qa_d,
      xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_21_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_21_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_21_i_1_inst_xt_rsc_0_21_i_qa_d_mxwt,
      xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_21_i_wea_d_pff => xt_rsc_0_21_i_wea_d_iff,
      xt_rsc_0_21_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_21_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_21_i_1_inst_xt_rsc_0_21_i_qa_d <= xt_rsc_0_21_i_qa_d;
  xt_rsc_0_21_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_21_i_1_inst_xt_rsc_0_21_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_22_i_1_inst : peaseNTT_core_xt_rsc_0_22_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_22_i_qa_d => peaseNTT_core_xt_rsc_0_22_i_1_inst_xt_rsc_0_22_i_qa_d,
      xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_22_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_22_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_22_i_1_inst_xt_rsc_0_22_i_qa_d_mxwt,
      xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_22_i_wea_d_pff => xt_rsc_0_22_i_wea_d_iff,
      xt_rsc_0_22_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_22_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_22_i_1_inst_xt_rsc_0_22_i_qa_d <= xt_rsc_0_22_i_qa_d;
  xt_rsc_0_22_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_22_i_1_inst_xt_rsc_0_22_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_23_i_1_inst : peaseNTT_core_xt_rsc_0_23_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_23_i_qa_d => peaseNTT_core_xt_rsc_0_23_i_1_inst_xt_rsc_0_23_i_qa_d,
      xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_23_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_23_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_23_i_1_inst_xt_rsc_0_23_i_qa_d_mxwt,
      xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_23_i_wea_d_pff => xt_rsc_0_23_i_wea_d_iff,
      xt_rsc_0_23_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_23_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_23_i_1_inst_xt_rsc_0_23_i_qa_d <= xt_rsc_0_23_i_qa_d;
  xt_rsc_0_23_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_23_i_1_inst_xt_rsc_0_23_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_24_i_1_inst : peaseNTT_core_xt_rsc_0_24_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_24_i_qa_d => peaseNTT_core_xt_rsc_0_24_i_1_inst_xt_rsc_0_24_i_qa_d,
      xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_24_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_24_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_24_i_1_inst_xt_rsc_0_24_i_qa_d_mxwt,
      xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_24_i_wea_d_pff => xt_rsc_0_24_i_wea_d_iff,
      xt_rsc_0_24_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_24_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_24_i_1_inst_xt_rsc_0_24_i_qa_d <= xt_rsc_0_24_i_qa_d;
  xt_rsc_0_24_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_24_i_1_inst_xt_rsc_0_24_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_25_i_1_inst : peaseNTT_core_xt_rsc_0_25_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_25_i_qa_d => peaseNTT_core_xt_rsc_0_25_i_1_inst_xt_rsc_0_25_i_qa_d,
      xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_25_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_25_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_25_i_1_inst_xt_rsc_0_25_i_qa_d_mxwt,
      xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_25_i_wea_d_pff => xt_rsc_0_25_i_wea_d_iff,
      xt_rsc_0_25_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_25_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_25_i_1_inst_xt_rsc_0_25_i_qa_d <= xt_rsc_0_25_i_qa_d;
  xt_rsc_0_25_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_25_i_1_inst_xt_rsc_0_25_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_26_i_1_inst : peaseNTT_core_xt_rsc_0_26_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_26_i_qa_d => peaseNTT_core_xt_rsc_0_26_i_1_inst_xt_rsc_0_26_i_qa_d,
      xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_26_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_26_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_26_i_1_inst_xt_rsc_0_26_i_qa_d_mxwt,
      xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_26_i_wea_d_pff => xt_rsc_0_26_i_wea_d_iff,
      xt_rsc_0_26_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_26_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_26_i_1_inst_xt_rsc_0_26_i_qa_d <= xt_rsc_0_26_i_qa_d;
  xt_rsc_0_26_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_26_i_1_inst_xt_rsc_0_26_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_27_i_1_inst : peaseNTT_core_xt_rsc_0_27_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_27_i_qa_d => peaseNTT_core_xt_rsc_0_27_i_1_inst_xt_rsc_0_27_i_qa_d,
      xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_27_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_27_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_27_i_1_inst_xt_rsc_0_27_i_qa_d_mxwt,
      xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_27_i_wea_d_pff => xt_rsc_0_27_i_wea_d_iff,
      xt_rsc_0_27_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_27_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_27_i_1_inst_xt_rsc_0_27_i_qa_d <= xt_rsc_0_27_i_qa_d;
  xt_rsc_0_27_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_27_i_1_inst_xt_rsc_0_27_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_28_i_1_inst : peaseNTT_core_xt_rsc_0_28_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_28_i_qa_d => peaseNTT_core_xt_rsc_0_28_i_1_inst_xt_rsc_0_28_i_qa_d,
      xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_28_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_28_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_28_i_1_inst_xt_rsc_0_28_i_qa_d_mxwt,
      xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_28_i_wea_d_pff => xt_rsc_0_28_i_wea_d_iff,
      xt_rsc_0_28_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_28_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_28_i_1_inst_xt_rsc_0_28_i_qa_d <= xt_rsc_0_28_i_qa_d;
  xt_rsc_0_28_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_28_i_1_inst_xt_rsc_0_28_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_29_i_1_inst : peaseNTT_core_xt_rsc_0_29_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_29_i_qa_d => peaseNTT_core_xt_rsc_0_29_i_1_inst_xt_rsc_0_29_i_qa_d,
      xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_29_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_29_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_29_i_1_inst_xt_rsc_0_29_i_qa_d_mxwt,
      xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_29_i_wea_d_pff => xt_rsc_0_29_i_wea_d_iff,
      xt_rsc_0_29_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_29_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_29_i_1_inst_xt_rsc_0_29_i_qa_d <= xt_rsc_0_29_i_qa_d;
  xt_rsc_0_29_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_29_i_1_inst_xt_rsc_0_29_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_30_i_1_inst : peaseNTT_core_xt_rsc_0_30_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_30_i_qa_d => peaseNTT_core_xt_rsc_0_30_i_1_inst_xt_rsc_0_30_i_qa_d,
      xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_30_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_30_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_30_i_1_inst_xt_rsc_0_30_i_qa_d_mxwt,
      xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_30_i_wea_d_pff => xt_rsc_0_30_i_wea_d_iff,
      xt_rsc_0_30_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_30_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_30_i_1_inst_xt_rsc_0_30_i_qa_d <= xt_rsc_0_30_i_qa_d;
  xt_rsc_0_30_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_30_i_1_inst_xt_rsc_0_30_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_0_31_i_1_inst : peaseNTT_core_xt_rsc_0_31_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_0_31_i_qa_d => peaseNTT_core_xt_rsc_0_31_i_1_inst_xt_rsc_0_31_i_qa_d,
      xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_0_31_i_oswt => reg_xt_rsc_0_16_i_oswt_cse,
      xt_rsc_0_31_i_qa_d_mxwt => peaseNTT_core_xt_rsc_0_31_i_1_inst_xt_rsc_0_31_i_qa_d_mxwt,
      xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_436_rmff,
      xt_rsc_0_31_i_wea_d_pff => xt_rsc_0_31_i_wea_d_iff,
      xt_rsc_0_31_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_0_31_i_oswt_pff => or_512_rmff
    );
  peaseNTT_core_xt_rsc_0_31_i_1_inst_xt_rsc_0_31_i_qa_d <= xt_rsc_0_31_i_qa_d;
  xt_rsc_0_31_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_0_31_i_1_inst_xt_rsc_0_31_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_0_i_1_inst : peaseNTT_core_xt_rsc_1_0_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_0_i_qa_d => peaseNTT_core_xt_rsc_1_0_i_1_inst_xt_rsc_1_0_i_qa_d,
      xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_0_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_0_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_0_i_1_inst_xt_rsc_1_0_i_qa_d_mxwt,
      xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_0_i_wea_d_pff => xt_rsc_1_0_i_wea_d_iff,
      xt_rsc_1_0_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_0_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_0_i_1_inst_xt_rsc_1_0_i_qa_d <= xt_rsc_1_0_i_qa_d;
  xt_rsc_1_0_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_0_i_1_inst_xt_rsc_1_0_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_1_i_1_inst : peaseNTT_core_xt_rsc_1_1_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_1_i_qa_d => peaseNTT_core_xt_rsc_1_1_i_1_inst_xt_rsc_1_1_i_qa_d,
      xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_1_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_1_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_1_i_1_inst_xt_rsc_1_1_i_qa_d_mxwt,
      xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_1_i_wea_d_pff => xt_rsc_1_1_i_wea_d_iff,
      xt_rsc_1_1_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_1_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_1_i_1_inst_xt_rsc_1_1_i_qa_d <= xt_rsc_1_1_i_qa_d;
  xt_rsc_1_1_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_1_i_1_inst_xt_rsc_1_1_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_2_i_1_inst : peaseNTT_core_xt_rsc_1_2_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_2_i_qa_d => peaseNTT_core_xt_rsc_1_2_i_1_inst_xt_rsc_1_2_i_qa_d,
      xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_2_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_2_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_2_i_1_inst_xt_rsc_1_2_i_qa_d_mxwt,
      xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_2_i_wea_d_pff => xt_rsc_1_2_i_wea_d_iff,
      xt_rsc_1_2_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_2_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_2_i_1_inst_xt_rsc_1_2_i_qa_d <= xt_rsc_1_2_i_qa_d;
  xt_rsc_1_2_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_2_i_1_inst_xt_rsc_1_2_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_3_i_1_inst : peaseNTT_core_xt_rsc_1_3_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_3_i_qa_d => peaseNTT_core_xt_rsc_1_3_i_1_inst_xt_rsc_1_3_i_qa_d,
      xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_3_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_3_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_3_i_1_inst_xt_rsc_1_3_i_qa_d_mxwt,
      xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_3_i_wea_d_pff => xt_rsc_1_3_i_wea_d_iff,
      xt_rsc_1_3_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_3_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_3_i_1_inst_xt_rsc_1_3_i_qa_d <= xt_rsc_1_3_i_qa_d;
  xt_rsc_1_3_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_3_i_1_inst_xt_rsc_1_3_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_4_i_1_inst : peaseNTT_core_xt_rsc_1_4_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_4_i_qa_d => peaseNTT_core_xt_rsc_1_4_i_1_inst_xt_rsc_1_4_i_qa_d,
      xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_4_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_4_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_4_i_1_inst_xt_rsc_1_4_i_qa_d_mxwt,
      xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_4_i_wea_d_pff => xt_rsc_1_4_i_wea_d_iff,
      xt_rsc_1_4_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_4_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_4_i_1_inst_xt_rsc_1_4_i_qa_d <= xt_rsc_1_4_i_qa_d;
  xt_rsc_1_4_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_4_i_1_inst_xt_rsc_1_4_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_5_i_1_inst : peaseNTT_core_xt_rsc_1_5_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_5_i_qa_d => peaseNTT_core_xt_rsc_1_5_i_1_inst_xt_rsc_1_5_i_qa_d,
      xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_5_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_5_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_5_i_1_inst_xt_rsc_1_5_i_qa_d_mxwt,
      xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_5_i_wea_d_pff => xt_rsc_1_5_i_wea_d_iff,
      xt_rsc_1_5_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_5_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_5_i_1_inst_xt_rsc_1_5_i_qa_d <= xt_rsc_1_5_i_qa_d;
  xt_rsc_1_5_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_5_i_1_inst_xt_rsc_1_5_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_6_i_1_inst : peaseNTT_core_xt_rsc_1_6_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_6_i_qa_d => peaseNTT_core_xt_rsc_1_6_i_1_inst_xt_rsc_1_6_i_qa_d,
      xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_6_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_6_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_6_i_1_inst_xt_rsc_1_6_i_qa_d_mxwt,
      xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_6_i_wea_d_pff => xt_rsc_1_6_i_wea_d_iff,
      xt_rsc_1_6_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_6_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_6_i_1_inst_xt_rsc_1_6_i_qa_d <= xt_rsc_1_6_i_qa_d;
  xt_rsc_1_6_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_6_i_1_inst_xt_rsc_1_6_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_7_i_1_inst : peaseNTT_core_xt_rsc_1_7_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_7_i_qa_d => peaseNTT_core_xt_rsc_1_7_i_1_inst_xt_rsc_1_7_i_qa_d,
      xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_7_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_7_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_7_i_1_inst_xt_rsc_1_7_i_qa_d_mxwt,
      xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_7_i_wea_d_pff => xt_rsc_1_7_i_wea_d_iff,
      xt_rsc_1_7_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_7_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_7_i_1_inst_xt_rsc_1_7_i_qa_d <= xt_rsc_1_7_i_qa_d;
  xt_rsc_1_7_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_7_i_1_inst_xt_rsc_1_7_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_8_i_1_inst : peaseNTT_core_xt_rsc_1_8_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_8_i_qa_d => peaseNTT_core_xt_rsc_1_8_i_1_inst_xt_rsc_1_8_i_qa_d,
      xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_8_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_8_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_8_i_1_inst_xt_rsc_1_8_i_qa_d_mxwt,
      xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_8_i_wea_d_pff => xt_rsc_1_8_i_wea_d_iff,
      xt_rsc_1_8_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_8_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_8_i_1_inst_xt_rsc_1_8_i_qa_d <= xt_rsc_1_8_i_qa_d;
  xt_rsc_1_8_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_8_i_1_inst_xt_rsc_1_8_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_9_i_1_inst : peaseNTT_core_xt_rsc_1_9_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_9_i_qa_d => peaseNTT_core_xt_rsc_1_9_i_1_inst_xt_rsc_1_9_i_qa_d,
      xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_9_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_9_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_9_i_1_inst_xt_rsc_1_9_i_qa_d_mxwt,
      xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_9_i_wea_d_pff => xt_rsc_1_9_i_wea_d_iff,
      xt_rsc_1_9_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_9_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_9_i_1_inst_xt_rsc_1_9_i_qa_d <= xt_rsc_1_9_i_qa_d;
  xt_rsc_1_9_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_9_i_1_inst_xt_rsc_1_9_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_10_i_1_inst : peaseNTT_core_xt_rsc_1_10_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_10_i_qa_d => peaseNTT_core_xt_rsc_1_10_i_1_inst_xt_rsc_1_10_i_qa_d,
      xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_10_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_10_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_10_i_1_inst_xt_rsc_1_10_i_qa_d_mxwt,
      xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_10_i_wea_d_pff => xt_rsc_1_10_i_wea_d_iff,
      xt_rsc_1_10_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_10_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_10_i_1_inst_xt_rsc_1_10_i_qa_d <= xt_rsc_1_10_i_qa_d;
  xt_rsc_1_10_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_10_i_1_inst_xt_rsc_1_10_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_11_i_1_inst : peaseNTT_core_xt_rsc_1_11_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_11_i_qa_d => peaseNTT_core_xt_rsc_1_11_i_1_inst_xt_rsc_1_11_i_qa_d,
      xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_11_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_11_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_11_i_1_inst_xt_rsc_1_11_i_qa_d_mxwt,
      xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_11_i_wea_d_pff => xt_rsc_1_11_i_wea_d_iff,
      xt_rsc_1_11_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_11_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_11_i_1_inst_xt_rsc_1_11_i_qa_d <= xt_rsc_1_11_i_qa_d;
  xt_rsc_1_11_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_11_i_1_inst_xt_rsc_1_11_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_12_i_1_inst : peaseNTT_core_xt_rsc_1_12_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_12_i_qa_d => peaseNTT_core_xt_rsc_1_12_i_1_inst_xt_rsc_1_12_i_qa_d,
      xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_12_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_12_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_12_i_1_inst_xt_rsc_1_12_i_qa_d_mxwt,
      xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_12_i_wea_d_pff => xt_rsc_1_12_i_wea_d_iff,
      xt_rsc_1_12_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_12_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_12_i_1_inst_xt_rsc_1_12_i_qa_d <= xt_rsc_1_12_i_qa_d;
  xt_rsc_1_12_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_12_i_1_inst_xt_rsc_1_12_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_13_i_1_inst : peaseNTT_core_xt_rsc_1_13_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_13_i_qa_d => peaseNTT_core_xt_rsc_1_13_i_1_inst_xt_rsc_1_13_i_qa_d,
      xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_13_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_13_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_13_i_1_inst_xt_rsc_1_13_i_qa_d_mxwt,
      xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_13_i_wea_d_pff => xt_rsc_1_13_i_wea_d_iff,
      xt_rsc_1_13_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_13_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_13_i_1_inst_xt_rsc_1_13_i_qa_d <= xt_rsc_1_13_i_qa_d;
  xt_rsc_1_13_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_13_i_1_inst_xt_rsc_1_13_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_14_i_1_inst : peaseNTT_core_xt_rsc_1_14_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_14_i_qa_d => peaseNTT_core_xt_rsc_1_14_i_1_inst_xt_rsc_1_14_i_qa_d,
      xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_14_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_14_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_14_i_1_inst_xt_rsc_1_14_i_qa_d_mxwt,
      xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_14_i_wea_d_pff => xt_rsc_1_14_i_wea_d_iff,
      xt_rsc_1_14_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_14_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_14_i_1_inst_xt_rsc_1_14_i_qa_d <= xt_rsc_1_14_i_qa_d;
  xt_rsc_1_14_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_14_i_1_inst_xt_rsc_1_14_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_15_i_1_inst : peaseNTT_core_xt_rsc_1_15_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_15_i_qa_d => peaseNTT_core_xt_rsc_1_15_i_1_inst_xt_rsc_1_15_i_qa_d,
      xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_15_i_oswt => reg_xt_rsc_1_0_i_oswt_cse,
      xt_rsc_1_15_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_15_i_1_inst_xt_rsc_1_15_i_qa_d_mxwt,
      xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_15_i_wea_d_pff => xt_rsc_1_15_i_wea_d_iff,
      xt_rsc_1_15_i_wea_d_core_psct_pff => or_435_rmff,
      xt_rsc_1_15_i_oswt_pff => or_578_rmff
    );
  peaseNTT_core_xt_rsc_1_15_i_1_inst_xt_rsc_1_15_i_qa_d <= xt_rsc_1_15_i_qa_d;
  xt_rsc_1_15_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_15_i_1_inst_xt_rsc_1_15_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_16_i_1_inst : peaseNTT_core_xt_rsc_1_16_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_16_i_qa_d => peaseNTT_core_xt_rsc_1_16_i_1_inst_xt_rsc_1_16_i_qa_d,
      xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_16_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_16_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_16_i_1_inst_xt_rsc_1_16_i_qa_d_mxwt,
      xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_16_i_wea_d_pff => xt_rsc_1_16_i_wea_d_iff,
      xt_rsc_1_16_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_16_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_16_i_1_inst_xt_rsc_1_16_i_qa_d <= xt_rsc_1_16_i_qa_d;
  xt_rsc_1_16_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_16_i_1_inst_xt_rsc_1_16_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_17_i_1_inst : peaseNTT_core_xt_rsc_1_17_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_17_i_qa_d => peaseNTT_core_xt_rsc_1_17_i_1_inst_xt_rsc_1_17_i_qa_d,
      xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_17_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_17_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_17_i_1_inst_xt_rsc_1_17_i_qa_d_mxwt,
      xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_17_i_wea_d_pff => xt_rsc_1_17_i_wea_d_iff,
      xt_rsc_1_17_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_17_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_17_i_1_inst_xt_rsc_1_17_i_qa_d <= xt_rsc_1_17_i_qa_d;
  xt_rsc_1_17_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_17_i_1_inst_xt_rsc_1_17_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_18_i_1_inst : peaseNTT_core_xt_rsc_1_18_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_18_i_qa_d => peaseNTT_core_xt_rsc_1_18_i_1_inst_xt_rsc_1_18_i_qa_d,
      xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_18_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_18_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_18_i_1_inst_xt_rsc_1_18_i_qa_d_mxwt,
      xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_18_i_wea_d_pff => xt_rsc_1_18_i_wea_d_iff,
      xt_rsc_1_18_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_18_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_18_i_1_inst_xt_rsc_1_18_i_qa_d <= xt_rsc_1_18_i_qa_d;
  xt_rsc_1_18_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_18_i_1_inst_xt_rsc_1_18_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_19_i_1_inst : peaseNTT_core_xt_rsc_1_19_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_19_i_qa_d => peaseNTT_core_xt_rsc_1_19_i_1_inst_xt_rsc_1_19_i_qa_d,
      xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_19_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_19_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_19_i_1_inst_xt_rsc_1_19_i_qa_d_mxwt,
      xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_19_i_wea_d_pff => xt_rsc_1_19_i_wea_d_iff,
      xt_rsc_1_19_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_19_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_19_i_1_inst_xt_rsc_1_19_i_qa_d <= xt_rsc_1_19_i_qa_d;
  xt_rsc_1_19_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_19_i_1_inst_xt_rsc_1_19_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_20_i_1_inst : peaseNTT_core_xt_rsc_1_20_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_20_i_qa_d => peaseNTT_core_xt_rsc_1_20_i_1_inst_xt_rsc_1_20_i_qa_d,
      xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_20_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_20_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_20_i_1_inst_xt_rsc_1_20_i_qa_d_mxwt,
      xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_20_i_wea_d_pff => xt_rsc_1_20_i_wea_d_iff,
      xt_rsc_1_20_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_20_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_20_i_1_inst_xt_rsc_1_20_i_qa_d <= xt_rsc_1_20_i_qa_d;
  xt_rsc_1_20_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_20_i_1_inst_xt_rsc_1_20_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_21_i_1_inst : peaseNTT_core_xt_rsc_1_21_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_21_i_qa_d => peaseNTT_core_xt_rsc_1_21_i_1_inst_xt_rsc_1_21_i_qa_d,
      xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_21_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_21_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_21_i_1_inst_xt_rsc_1_21_i_qa_d_mxwt,
      xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_21_i_wea_d_pff => xt_rsc_1_21_i_wea_d_iff,
      xt_rsc_1_21_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_21_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_21_i_1_inst_xt_rsc_1_21_i_qa_d <= xt_rsc_1_21_i_qa_d;
  xt_rsc_1_21_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_21_i_1_inst_xt_rsc_1_21_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_22_i_1_inst : peaseNTT_core_xt_rsc_1_22_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_22_i_qa_d => peaseNTT_core_xt_rsc_1_22_i_1_inst_xt_rsc_1_22_i_qa_d,
      xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_22_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_22_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_22_i_1_inst_xt_rsc_1_22_i_qa_d_mxwt,
      xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_22_i_wea_d_pff => xt_rsc_1_22_i_wea_d_iff,
      xt_rsc_1_22_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_22_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_22_i_1_inst_xt_rsc_1_22_i_qa_d <= xt_rsc_1_22_i_qa_d;
  xt_rsc_1_22_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_22_i_1_inst_xt_rsc_1_22_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_23_i_1_inst : peaseNTT_core_xt_rsc_1_23_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_23_i_qa_d => peaseNTT_core_xt_rsc_1_23_i_1_inst_xt_rsc_1_23_i_qa_d,
      xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_23_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_23_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_23_i_1_inst_xt_rsc_1_23_i_qa_d_mxwt,
      xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_23_i_wea_d_pff => xt_rsc_1_23_i_wea_d_iff,
      xt_rsc_1_23_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_23_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_23_i_1_inst_xt_rsc_1_23_i_qa_d <= xt_rsc_1_23_i_qa_d;
  xt_rsc_1_23_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_23_i_1_inst_xt_rsc_1_23_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_24_i_1_inst : peaseNTT_core_xt_rsc_1_24_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_24_i_qa_d => peaseNTT_core_xt_rsc_1_24_i_1_inst_xt_rsc_1_24_i_qa_d,
      xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_24_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_24_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_24_i_1_inst_xt_rsc_1_24_i_qa_d_mxwt,
      xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_24_i_wea_d_pff => xt_rsc_1_24_i_wea_d_iff,
      xt_rsc_1_24_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_24_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_24_i_1_inst_xt_rsc_1_24_i_qa_d <= xt_rsc_1_24_i_qa_d;
  xt_rsc_1_24_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_24_i_1_inst_xt_rsc_1_24_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_25_i_1_inst : peaseNTT_core_xt_rsc_1_25_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_25_i_qa_d => peaseNTT_core_xt_rsc_1_25_i_1_inst_xt_rsc_1_25_i_qa_d,
      xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_25_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_25_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_25_i_1_inst_xt_rsc_1_25_i_qa_d_mxwt,
      xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_25_i_wea_d_pff => xt_rsc_1_25_i_wea_d_iff,
      xt_rsc_1_25_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_25_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_25_i_1_inst_xt_rsc_1_25_i_qa_d <= xt_rsc_1_25_i_qa_d;
  xt_rsc_1_25_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_25_i_1_inst_xt_rsc_1_25_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_26_i_1_inst : peaseNTT_core_xt_rsc_1_26_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_26_i_qa_d => peaseNTT_core_xt_rsc_1_26_i_1_inst_xt_rsc_1_26_i_qa_d,
      xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_26_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_26_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_26_i_1_inst_xt_rsc_1_26_i_qa_d_mxwt,
      xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_26_i_wea_d_pff => xt_rsc_1_26_i_wea_d_iff,
      xt_rsc_1_26_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_26_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_26_i_1_inst_xt_rsc_1_26_i_qa_d <= xt_rsc_1_26_i_qa_d;
  xt_rsc_1_26_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_26_i_1_inst_xt_rsc_1_26_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_27_i_1_inst : peaseNTT_core_xt_rsc_1_27_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_27_i_qa_d => peaseNTT_core_xt_rsc_1_27_i_1_inst_xt_rsc_1_27_i_qa_d,
      xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_27_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_27_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_27_i_1_inst_xt_rsc_1_27_i_qa_d_mxwt,
      xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_27_i_wea_d_pff => xt_rsc_1_27_i_wea_d_iff,
      xt_rsc_1_27_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_27_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_27_i_1_inst_xt_rsc_1_27_i_qa_d <= xt_rsc_1_27_i_qa_d;
  xt_rsc_1_27_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_27_i_1_inst_xt_rsc_1_27_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_28_i_1_inst : peaseNTT_core_xt_rsc_1_28_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_28_i_qa_d => peaseNTT_core_xt_rsc_1_28_i_1_inst_xt_rsc_1_28_i_qa_d,
      xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_28_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_28_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_28_i_1_inst_xt_rsc_1_28_i_qa_d_mxwt,
      xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_28_i_wea_d_pff => xt_rsc_1_28_i_wea_d_iff,
      xt_rsc_1_28_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_28_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_28_i_1_inst_xt_rsc_1_28_i_qa_d <= xt_rsc_1_28_i_qa_d;
  xt_rsc_1_28_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_28_i_1_inst_xt_rsc_1_28_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_29_i_1_inst : peaseNTT_core_xt_rsc_1_29_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_29_i_qa_d => peaseNTT_core_xt_rsc_1_29_i_1_inst_xt_rsc_1_29_i_qa_d,
      xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_29_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_29_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_29_i_1_inst_xt_rsc_1_29_i_qa_d_mxwt,
      xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_29_i_wea_d_pff => xt_rsc_1_29_i_wea_d_iff,
      xt_rsc_1_29_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_29_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_29_i_1_inst_xt_rsc_1_29_i_qa_d <= xt_rsc_1_29_i_qa_d;
  xt_rsc_1_29_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_29_i_1_inst_xt_rsc_1_29_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_30_i_1_inst : peaseNTT_core_xt_rsc_1_30_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_30_i_qa_d => peaseNTT_core_xt_rsc_1_30_i_1_inst_xt_rsc_1_30_i_qa_d,
      xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_30_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_30_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_30_i_1_inst_xt_rsc_1_30_i_qa_d_mxwt,
      xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_30_i_wea_d_pff => xt_rsc_1_30_i_wea_d_iff,
      xt_rsc_1_30_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_30_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_30_i_1_inst_xt_rsc_1_30_i_qa_d <= xt_rsc_1_30_i_qa_d;
  xt_rsc_1_30_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_30_i_1_inst_xt_rsc_1_30_i_qa_d_mxwt;

  peaseNTT_core_xt_rsc_1_31_i_1_inst : peaseNTT_core_xt_rsc_1_31_i_1
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_1_31_i_qa_d => peaseNTT_core_xt_rsc_1_31_i_1_inst_xt_rsc_1_31_i_qa_d,
      xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg,
      core_wen => core_wen,
      core_wten => core_wten,
      xt_rsc_1_31_i_oswt => reg_xt_rsc_1_16_i_oswt_cse,
      xt_rsc_1_31_i_qa_d_mxwt => peaseNTT_core_xt_rsc_1_31_i_1_inst_xt_rsc_1_31_i_qa_d_mxwt,
      xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_core_psct => or_584_rmff,
      xt_rsc_1_31_i_wea_d_pff => xt_rsc_1_31_i_wea_d_iff,
      xt_rsc_1_31_i_wea_d_core_psct_pff => or_517_rmff,
      xt_rsc_1_31_i_oswt_pff => or_660_rmff
    );
  peaseNTT_core_xt_rsc_1_31_i_1_inst_xt_rsc_1_31_i_qa_d <= xt_rsc_1_31_i_qa_d;
  xt_rsc_1_31_i_qa_d_mxwt <= peaseNTT_core_xt_rsc_1_31_i_1_inst_xt_rsc_1_31_i_qa_d_mxwt;

  peaseNTT_core_twiddle_rsc_0_0_i_inst : peaseNTT_core_twiddle_rsc_0_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_0_s_tdone => twiddle_rsc_0_0_s_tdone,
      twiddle_rsc_0_0_tr_write_done => twiddle_rsc_0_0_tr_write_done,
      twiddle_rsc_0_0_RREADY => twiddle_rsc_0_0_RREADY,
      twiddle_rsc_0_0_RVALID => twiddle_rsc_0_0_RVALID,
      twiddle_rsc_0_0_RUSER => twiddle_rsc_0_0_RUSER,
      twiddle_rsc_0_0_RLAST => twiddle_rsc_0_0_RLAST,
      twiddle_rsc_0_0_RRESP => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_RRESP,
      twiddle_rsc_0_0_RDATA => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_RDATA,
      twiddle_rsc_0_0_RID => twiddle_rsc_0_0_RID,
      twiddle_rsc_0_0_ARREADY => twiddle_rsc_0_0_ARREADY,
      twiddle_rsc_0_0_ARVALID => twiddle_rsc_0_0_ARVALID,
      twiddle_rsc_0_0_ARUSER => twiddle_rsc_0_0_ARUSER,
      twiddle_rsc_0_0_ARREGION => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARREGION,
      twiddle_rsc_0_0_ARQOS => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARQOS,
      twiddle_rsc_0_0_ARPROT => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARPROT,
      twiddle_rsc_0_0_ARCACHE => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARCACHE,
      twiddle_rsc_0_0_ARLOCK => twiddle_rsc_0_0_ARLOCK,
      twiddle_rsc_0_0_ARBURST => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARBURST,
      twiddle_rsc_0_0_ARSIZE => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARSIZE,
      twiddle_rsc_0_0_ARLEN => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARLEN,
      twiddle_rsc_0_0_ARADDR => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARADDR,
      twiddle_rsc_0_0_ARID => twiddle_rsc_0_0_ARID,
      twiddle_rsc_0_0_BREADY => twiddle_rsc_0_0_BREADY,
      twiddle_rsc_0_0_BVALID => twiddle_rsc_0_0_BVALID,
      twiddle_rsc_0_0_BUSER => twiddle_rsc_0_0_BUSER,
      twiddle_rsc_0_0_BRESP => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_BRESP,
      twiddle_rsc_0_0_BID => twiddle_rsc_0_0_BID,
      twiddle_rsc_0_0_WREADY => twiddle_rsc_0_0_WREADY,
      twiddle_rsc_0_0_WVALID => twiddle_rsc_0_0_WVALID,
      twiddle_rsc_0_0_WUSER => twiddle_rsc_0_0_WUSER,
      twiddle_rsc_0_0_WLAST => twiddle_rsc_0_0_WLAST,
      twiddle_rsc_0_0_WSTRB => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_WSTRB,
      twiddle_rsc_0_0_WDATA => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_WDATA,
      twiddle_rsc_0_0_AWREADY => twiddle_rsc_0_0_AWREADY,
      twiddle_rsc_0_0_AWVALID => twiddle_rsc_0_0_AWVALID,
      twiddle_rsc_0_0_AWUSER => twiddle_rsc_0_0_AWUSER,
      twiddle_rsc_0_0_AWREGION => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWREGION,
      twiddle_rsc_0_0_AWQOS => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWQOS,
      twiddle_rsc_0_0_AWPROT => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWPROT,
      twiddle_rsc_0_0_AWCACHE => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWCACHE,
      twiddle_rsc_0_0_AWLOCK => twiddle_rsc_0_0_AWLOCK,
      twiddle_rsc_0_0_AWBURST => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWBURST,
      twiddle_rsc_0_0_AWSIZE => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWSIZE,
      twiddle_rsc_0_0_AWLEN => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWLEN,
      twiddle_rsc_0_0_AWADDR => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWADDR,
      twiddle_rsc_0_0_AWID => twiddle_rsc_0_0_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_0_i_oswt => reg_twiddle_rsc_0_0_i_oswt_cse,
      twiddle_rsc_0_0_i_wen_comp => twiddle_rsc_0_0_i_wen_comp,
      twiddle_rsc_0_0_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_i_s_raddr_core,
      twiddle_rsc_0_0_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_i_s_din_mxwt
    );
  twiddle_rsc_0_0_RRESP <= peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_RRESP;
  twiddle_rsc_0_0_RDATA <= peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_RDATA;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARREGION <= twiddle_rsc_0_0_ARREGION;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARQOS <= twiddle_rsc_0_0_ARQOS;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARPROT <= twiddle_rsc_0_0_ARPROT;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARCACHE <= twiddle_rsc_0_0_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARBURST <= twiddle_rsc_0_0_ARBURST;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARSIZE <= twiddle_rsc_0_0_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARLEN <= twiddle_rsc_0_0_ARLEN;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_ARADDR <= twiddle_rsc_0_0_ARADDR;
  twiddle_rsc_0_0_BRESP <= peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_BRESP;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_WSTRB <= twiddle_rsc_0_0_WSTRB;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_WDATA <= twiddle_rsc_0_0_WDATA;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWREGION <= twiddle_rsc_0_0_AWREGION;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWQOS <= twiddle_rsc_0_0_AWQOS;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWPROT <= twiddle_rsc_0_0_AWPROT;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWCACHE <= twiddle_rsc_0_0_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWBURST <= twiddle_rsc_0_0_AWBURST;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWSIZE <= twiddle_rsc_0_0_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWLEN <= twiddle_rsc_0_0_AWLEN;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_AWADDR <= twiddle_rsc_0_0_AWADDR;
  peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_i_s_raddr_core <= '0' & twiddle_h_rsc_0_0_i_s_raddr_core_4
      & reg_twiddle_rsc_0_0_i_s_raddr_core_3_0_cse;
  twiddle_rsc_0_0_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_0_i_inst_twiddle_rsc_0_0_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_1_i_inst : peaseNTT_core_twiddle_rsc_0_1_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_1_s_tdone => twiddle_rsc_0_1_s_tdone,
      twiddle_rsc_0_1_tr_write_done => twiddle_rsc_0_1_tr_write_done,
      twiddle_rsc_0_1_RREADY => twiddle_rsc_0_1_RREADY,
      twiddle_rsc_0_1_RVALID => twiddle_rsc_0_1_RVALID,
      twiddle_rsc_0_1_RUSER => twiddle_rsc_0_1_RUSER,
      twiddle_rsc_0_1_RLAST => twiddle_rsc_0_1_RLAST,
      twiddle_rsc_0_1_RRESP => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_RRESP,
      twiddle_rsc_0_1_RDATA => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_RDATA,
      twiddle_rsc_0_1_RID => twiddle_rsc_0_1_RID,
      twiddle_rsc_0_1_ARREADY => twiddle_rsc_0_1_ARREADY,
      twiddle_rsc_0_1_ARVALID => twiddle_rsc_0_1_ARVALID,
      twiddle_rsc_0_1_ARUSER => twiddle_rsc_0_1_ARUSER,
      twiddle_rsc_0_1_ARREGION => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARREGION,
      twiddle_rsc_0_1_ARQOS => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARQOS,
      twiddle_rsc_0_1_ARPROT => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARPROT,
      twiddle_rsc_0_1_ARCACHE => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARCACHE,
      twiddle_rsc_0_1_ARLOCK => twiddle_rsc_0_1_ARLOCK,
      twiddle_rsc_0_1_ARBURST => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARBURST,
      twiddle_rsc_0_1_ARSIZE => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARSIZE,
      twiddle_rsc_0_1_ARLEN => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARLEN,
      twiddle_rsc_0_1_ARADDR => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARADDR,
      twiddle_rsc_0_1_ARID => twiddle_rsc_0_1_ARID,
      twiddle_rsc_0_1_BREADY => twiddle_rsc_0_1_BREADY,
      twiddle_rsc_0_1_BVALID => twiddle_rsc_0_1_BVALID,
      twiddle_rsc_0_1_BUSER => twiddle_rsc_0_1_BUSER,
      twiddle_rsc_0_1_BRESP => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_BRESP,
      twiddle_rsc_0_1_BID => twiddle_rsc_0_1_BID,
      twiddle_rsc_0_1_WREADY => twiddle_rsc_0_1_WREADY,
      twiddle_rsc_0_1_WVALID => twiddle_rsc_0_1_WVALID,
      twiddle_rsc_0_1_WUSER => twiddle_rsc_0_1_WUSER,
      twiddle_rsc_0_1_WLAST => twiddle_rsc_0_1_WLAST,
      twiddle_rsc_0_1_WSTRB => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_WSTRB,
      twiddle_rsc_0_1_WDATA => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_WDATA,
      twiddle_rsc_0_1_AWREADY => twiddle_rsc_0_1_AWREADY,
      twiddle_rsc_0_1_AWVALID => twiddle_rsc_0_1_AWVALID,
      twiddle_rsc_0_1_AWUSER => twiddle_rsc_0_1_AWUSER,
      twiddle_rsc_0_1_AWREGION => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWREGION,
      twiddle_rsc_0_1_AWQOS => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWQOS,
      twiddle_rsc_0_1_AWPROT => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWPROT,
      twiddle_rsc_0_1_AWCACHE => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWCACHE,
      twiddle_rsc_0_1_AWLOCK => twiddle_rsc_0_1_AWLOCK,
      twiddle_rsc_0_1_AWBURST => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWBURST,
      twiddle_rsc_0_1_AWSIZE => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWSIZE,
      twiddle_rsc_0_1_AWLEN => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWLEN,
      twiddle_rsc_0_1_AWADDR => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWADDR,
      twiddle_rsc_0_1_AWID => twiddle_rsc_0_1_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_1_i_oswt => reg_twiddle_rsc_0_1_i_oswt_cse,
      twiddle_rsc_0_1_i_wen_comp => twiddle_rsc_0_1_i_wen_comp,
      twiddle_rsc_0_1_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_i_s_raddr_core,
      twiddle_rsc_0_1_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_i_s_din_mxwt
    );
  twiddle_rsc_0_1_RRESP <= peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_RRESP;
  twiddle_rsc_0_1_RDATA <= peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_RDATA;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARREGION <= twiddle_rsc_0_1_ARREGION;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARQOS <= twiddle_rsc_0_1_ARQOS;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARPROT <= twiddle_rsc_0_1_ARPROT;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARCACHE <= twiddle_rsc_0_1_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARBURST <= twiddle_rsc_0_1_ARBURST;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARSIZE <= twiddle_rsc_0_1_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARLEN <= twiddle_rsc_0_1_ARLEN;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_ARADDR <= twiddle_rsc_0_1_ARADDR;
  twiddle_rsc_0_1_BRESP <= peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_BRESP;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_WSTRB <= twiddle_rsc_0_1_WSTRB;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_WDATA <= twiddle_rsc_0_1_WDATA;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWREGION <= twiddle_rsc_0_1_AWREGION;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWQOS <= twiddle_rsc_0_1_AWQOS;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWPROT <= twiddle_rsc_0_1_AWPROT;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWCACHE <= twiddle_rsc_0_1_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWBURST <= twiddle_rsc_0_1_AWBURST;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWSIZE <= twiddle_rsc_0_1_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWLEN <= twiddle_rsc_0_1_AWLEN;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_AWADDR <= twiddle_rsc_0_1_AWADDR;
  peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_1_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_1_i_inst_twiddle_rsc_0_1_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_2_i_inst : peaseNTT_core_twiddle_rsc_0_2_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_2_s_tdone => twiddle_rsc_0_2_s_tdone,
      twiddle_rsc_0_2_tr_write_done => twiddle_rsc_0_2_tr_write_done,
      twiddle_rsc_0_2_RREADY => twiddle_rsc_0_2_RREADY,
      twiddle_rsc_0_2_RVALID => twiddle_rsc_0_2_RVALID,
      twiddle_rsc_0_2_RUSER => twiddle_rsc_0_2_RUSER,
      twiddle_rsc_0_2_RLAST => twiddle_rsc_0_2_RLAST,
      twiddle_rsc_0_2_RRESP => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_RRESP,
      twiddle_rsc_0_2_RDATA => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_RDATA,
      twiddle_rsc_0_2_RID => twiddle_rsc_0_2_RID,
      twiddle_rsc_0_2_ARREADY => twiddle_rsc_0_2_ARREADY,
      twiddle_rsc_0_2_ARVALID => twiddle_rsc_0_2_ARVALID,
      twiddle_rsc_0_2_ARUSER => twiddle_rsc_0_2_ARUSER,
      twiddle_rsc_0_2_ARREGION => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARREGION,
      twiddle_rsc_0_2_ARQOS => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARQOS,
      twiddle_rsc_0_2_ARPROT => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARPROT,
      twiddle_rsc_0_2_ARCACHE => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARCACHE,
      twiddle_rsc_0_2_ARLOCK => twiddle_rsc_0_2_ARLOCK,
      twiddle_rsc_0_2_ARBURST => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARBURST,
      twiddle_rsc_0_2_ARSIZE => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARSIZE,
      twiddle_rsc_0_2_ARLEN => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARLEN,
      twiddle_rsc_0_2_ARADDR => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARADDR,
      twiddle_rsc_0_2_ARID => twiddle_rsc_0_2_ARID,
      twiddle_rsc_0_2_BREADY => twiddle_rsc_0_2_BREADY,
      twiddle_rsc_0_2_BVALID => twiddle_rsc_0_2_BVALID,
      twiddle_rsc_0_2_BUSER => twiddle_rsc_0_2_BUSER,
      twiddle_rsc_0_2_BRESP => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_BRESP,
      twiddle_rsc_0_2_BID => twiddle_rsc_0_2_BID,
      twiddle_rsc_0_2_WREADY => twiddle_rsc_0_2_WREADY,
      twiddle_rsc_0_2_WVALID => twiddle_rsc_0_2_WVALID,
      twiddle_rsc_0_2_WUSER => twiddle_rsc_0_2_WUSER,
      twiddle_rsc_0_2_WLAST => twiddle_rsc_0_2_WLAST,
      twiddle_rsc_0_2_WSTRB => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_WSTRB,
      twiddle_rsc_0_2_WDATA => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_WDATA,
      twiddle_rsc_0_2_AWREADY => twiddle_rsc_0_2_AWREADY,
      twiddle_rsc_0_2_AWVALID => twiddle_rsc_0_2_AWVALID,
      twiddle_rsc_0_2_AWUSER => twiddle_rsc_0_2_AWUSER,
      twiddle_rsc_0_2_AWREGION => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWREGION,
      twiddle_rsc_0_2_AWQOS => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWQOS,
      twiddle_rsc_0_2_AWPROT => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWPROT,
      twiddle_rsc_0_2_AWCACHE => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWCACHE,
      twiddle_rsc_0_2_AWLOCK => twiddle_rsc_0_2_AWLOCK,
      twiddle_rsc_0_2_AWBURST => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWBURST,
      twiddle_rsc_0_2_AWSIZE => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWSIZE,
      twiddle_rsc_0_2_AWLEN => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWLEN,
      twiddle_rsc_0_2_AWADDR => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWADDR,
      twiddle_rsc_0_2_AWID => twiddle_rsc_0_2_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_2_i_oswt => reg_twiddle_rsc_0_2_i_oswt_cse,
      twiddle_rsc_0_2_i_wen_comp => twiddle_rsc_0_2_i_wen_comp,
      twiddle_rsc_0_2_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_i_s_raddr_core,
      twiddle_rsc_0_2_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_i_s_din_mxwt
    );
  twiddle_rsc_0_2_RRESP <= peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_RRESP;
  twiddle_rsc_0_2_RDATA <= peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_RDATA;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARREGION <= twiddle_rsc_0_2_ARREGION;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARQOS <= twiddle_rsc_0_2_ARQOS;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARPROT <= twiddle_rsc_0_2_ARPROT;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARCACHE <= twiddle_rsc_0_2_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARBURST <= twiddle_rsc_0_2_ARBURST;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARSIZE <= twiddle_rsc_0_2_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARLEN <= twiddle_rsc_0_2_ARLEN;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_ARADDR <= twiddle_rsc_0_2_ARADDR;
  twiddle_rsc_0_2_BRESP <= peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_BRESP;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_WSTRB <= twiddle_rsc_0_2_WSTRB;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_WDATA <= twiddle_rsc_0_2_WDATA;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWREGION <= twiddle_rsc_0_2_AWREGION;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWQOS <= twiddle_rsc_0_2_AWQOS;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWPROT <= twiddle_rsc_0_2_AWPROT;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWCACHE <= twiddle_rsc_0_2_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWBURST <= twiddle_rsc_0_2_AWBURST;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWSIZE <= twiddle_rsc_0_2_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWLEN <= twiddle_rsc_0_2_AWLEN;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_AWADDR <= twiddle_rsc_0_2_AWADDR;
  peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_2_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_2_i_inst_twiddle_rsc_0_2_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_3_i_inst : peaseNTT_core_twiddle_rsc_0_3_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_3_s_tdone => twiddle_rsc_0_3_s_tdone,
      twiddle_rsc_0_3_tr_write_done => twiddle_rsc_0_3_tr_write_done,
      twiddle_rsc_0_3_RREADY => twiddle_rsc_0_3_RREADY,
      twiddle_rsc_0_3_RVALID => twiddle_rsc_0_3_RVALID,
      twiddle_rsc_0_3_RUSER => twiddle_rsc_0_3_RUSER,
      twiddle_rsc_0_3_RLAST => twiddle_rsc_0_3_RLAST,
      twiddle_rsc_0_3_RRESP => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_RRESP,
      twiddle_rsc_0_3_RDATA => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_RDATA,
      twiddle_rsc_0_3_RID => twiddle_rsc_0_3_RID,
      twiddle_rsc_0_3_ARREADY => twiddle_rsc_0_3_ARREADY,
      twiddle_rsc_0_3_ARVALID => twiddle_rsc_0_3_ARVALID,
      twiddle_rsc_0_3_ARUSER => twiddle_rsc_0_3_ARUSER,
      twiddle_rsc_0_3_ARREGION => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARREGION,
      twiddle_rsc_0_3_ARQOS => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARQOS,
      twiddle_rsc_0_3_ARPROT => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARPROT,
      twiddle_rsc_0_3_ARCACHE => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARCACHE,
      twiddle_rsc_0_3_ARLOCK => twiddle_rsc_0_3_ARLOCK,
      twiddle_rsc_0_3_ARBURST => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARBURST,
      twiddle_rsc_0_3_ARSIZE => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARSIZE,
      twiddle_rsc_0_3_ARLEN => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARLEN,
      twiddle_rsc_0_3_ARADDR => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARADDR,
      twiddle_rsc_0_3_ARID => twiddle_rsc_0_3_ARID,
      twiddle_rsc_0_3_BREADY => twiddle_rsc_0_3_BREADY,
      twiddle_rsc_0_3_BVALID => twiddle_rsc_0_3_BVALID,
      twiddle_rsc_0_3_BUSER => twiddle_rsc_0_3_BUSER,
      twiddle_rsc_0_3_BRESP => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_BRESP,
      twiddle_rsc_0_3_BID => twiddle_rsc_0_3_BID,
      twiddle_rsc_0_3_WREADY => twiddle_rsc_0_3_WREADY,
      twiddle_rsc_0_3_WVALID => twiddle_rsc_0_3_WVALID,
      twiddle_rsc_0_3_WUSER => twiddle_rsc_0_3_WUSER,
      twiddle_rsc_0_3_WLAST => twiddle_rsc_0_3_WLAST,
      twiddle_rsc_0_3_WSTRB => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_WSTRB,
      twiddle_rsc_0_3_WDATA => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_WDATA,
      twiddle_rsc_0_3_AWREADY => twiddle_rsc_0_3_AWREADY,
      twiddle_rsc_0_3_AWVALID => twiddle_rsc_0_3_AWVALID,
      twiddle_rsc_0_3_AWUSER => twiddle_rsc_0_3_AWUSER,
      twiddle_rsc_0_3_AWREGION => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWREGION,
      twiddle_rsc_0_3_AWQOS => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWQOS,
      twiddle_rsc_0_3_AWPROT => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWPROT,
      twiddle_rsc_0_3_AWCACHE => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWCACHE,
      twiddle_rsc_0_3_AWLOCK => twiddle_rsc_0_3_AWLOCK,
      twiddle_rsc_0_3_AWBURST => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWBURST,
      twiddle_rsc_0_3_AWSIZE => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWSIZE,
      twiddle_rsc_0_3_AWLEN => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWLEN,
      twiddle_rsc_0_3_AWADDR => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWADDR,
      twiddle_rsc_0_3_AWID => twiddle_rsc_0_3_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_3_i_oswt => reg_twiddle_rsc_0_3_i_oswt_cse,
      twiddle_rsc_0_3_i_wen_comp => twiddle_rsc_0_3_i_wen_comp,
      twiddle_rsc_0_3_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_i_s_raddr_core,
      twiddle_rsc_0_3_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_i_s_din_mxwt
    );
  twiddle_rsc_0_3_RRESP <= peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_RRESP;
  twiddle_rsc_0_3_RDATA <= peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_RDATA;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARREGION <= twiddle_rsc_0_3_ARREGION;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARQOS <= twiddle_rsc_0_3_ARQOS;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARPROT <= twiddle_rsc_0_3_ARPROT;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARCACHE <= twiddle_rsc_0_3_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARBURST <= twiddle_rsc_0_3_ARBURST;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARSIZE <= twiddle_rsc_0_3_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARLEN <= twiddle_rsc_0_3_ARLEN;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_ARADDR <= twiddle_rsc_0_3_ARADDR;
  twiddle_rsc_0_3_BRESP <= peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_BRESP;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_WSTRB <= twiddle_rsc_0_3_WSTRB;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_WDATA <= twiddle_rsc_0_3_WDATA;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWREGION <= twiddle_rsc_0_3_AWREGION;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWQOS <= twiddle_rsc_0_3_AWQOS;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWPROT <= twiddle_rsc_0_3_AWPROT;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWCACHE <= twiddle_rsc_0_3_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWBURST <= twiddle_rsc_0_3_AWBURST;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWSIZE <= twiddle_rsc_0_3_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWLEN <= twiddle_rsc_0_3_AWLEN;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_AWADDR <= twiddle_rsc_0_3_AWADDR;
  peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_3_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_3_i_inst_twiddle_rsc_0_3_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_4_i_inst : peaseNTT_core_twiddle_rsc_0_4_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_4_s_tdone => twiddle_rsc_0_4_s_tdone,
      twiddle_rsc_0_4_tr_write_done => twiddle_rsc_0_4_tr_write_done,
      twiddle_rsc_0_4_RREADY => twiddle_rsc_0_4_RREADY,
      twiddle_rsc_0_4_RVALID => twiddle_rsc_0_4_RVALID,
      twiddle_rsc_0_4_RUSER => twiddle_rsc_0_4_RUSER,
      twiddle_rsc_0_4_RLAST => twiddle_rsc_0_4_RLAST,
      twiddle_rsc_0_4_RRESP => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_RRESP,
      twiddle_rsc_0_4_RDATA => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_RDATA,
      twiddle_rsc_0_4_RID => twiddle_rsc_0_4_RID,
      twiddle_rsc_0_4_ARREADY => twiddle_rsc_0_4_ARREADY,
      twiddle_rsc_0_4_ARVALID => twiddle_rsc_0_4_ARVALID,
      twiddle_rsc_0_4_ARUSER => twiddle_rsc_0_4_ARUSER,
      twiddle_rsc_0_4_ARREGION => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARREGION,
      twiddle_rsc_0_4_ARQOS => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARQOS,
      twiddle_rsc_0_4_ARPROT => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARPROT,
      twiddle_rsc_0_4_ARCACHE => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARCACHE,
      twiddle_rsc_0_4_ARLOCK => twiddle_rsc_0_4_ARLOCK,
      twiddle_rsc_0_4_ARBURST => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARBURST,
      twiddle_rsc_0_4_ARSIZE => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARSIZE,
      twiddle_rsc_0_4_ARLEN => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARLEN,
      twiddle_rsc_0_4_ARADDR => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARADDR,
      twiddle_rsc_0_4_ARID => twiddle_rsc_0_4_ARID,
      twiddle_rsc_0_4_BREADY => twiddle_rsc_0_4_BREADY,
      twiddle_rsc_0_4_BVALID => twiddle_rsc_0_4_BVALID,
      twiddle_rsc_0_4_BUSER => twiddle_rsc_0_4_BUSER,
      twiddle_rsc_0_4_BRESP => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_BRESP,
      twiddle_rsc_0_4_BID => twiddle_rsc_0_4_BID,
      twiddle_rsc_0_4_WREADY => twiddle_rsc_0_4_WREADY,
      twiddle_rsc_0_4_WVALID => twiddle_rsc_0_4_WVALID,
      twiddle_rsc_0_4_WUSER => twiddle_rsc_0_4_WUSER,
      twiddle_rsc_0_4_WLAST => twiddle_rsc_0_4_WLAST,
      twiddle_rsc_0_4_WSTRB => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_WSTRB,
      twiddle_rsc_0_4_WDATA => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_WDATA,
      twiddle_rsc_0_4_AWREADY => twiddle_rsc_0_4_AWREADY,
      twiddle_rsc_0_4_AWVALID => twiddle_rsc_0_4_AWVALID,
      twiddle_rsc_0_4_AWUSER => twiddle_rsc_0_4_AWUSER,
      twiddle_rsc_0_4_AWREGION => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWREGION,
      twiddle_rsc_0_4_AWQOS => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWQOS,
      twiddle_rsc_0_4_AWPROT => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWPROT,
      twiddle_rsc_0_4_AWCACHE => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWCACHE,
      twiddle_rsc_0_4_AWLOCK => twiddle_rsc_0_4_AWLOCK,
      twiddle_rsc_0_4_AWBURST => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWBURST,
      twiddle_rsc_0_4_AWSIZE => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWSIZE,
      twiddle_rsc_0_4_AWLEN => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWLEN,
      twiddle_rsc_0_4_AWADDR => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWADDR,
      twiddle_rsc_0_4_AWID => twiddle_rsc_0_4_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_4_i_oswt => reg_twiddle_rsc_0_4_i_oswt_cse,
      twiddle_rsc_0_4_i_wen_comp => twiddle_rsc_0_4_i_wen_comp,
      twiddle_rsc_0_4_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_i_s_raddr_core,
      twiddle_rsc_0_4_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_i_s_din_mxwt
    );
  twiddle_rsc_0_4_RRESP <= peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_RRESP;
  twiddle_rsc_0_4_RDATA <= peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_RDATA;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARREGION <= twiddle_rsc_0_4_ARREGION;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARQOS <= twiddle_rsc_0_4_ARQOS;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARPROT <= twiddle_rsc_0_4_ARPROT;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARCACHE <= twiddle_rsc_0_4_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARBURST <= twiddle_rsc_0_4_ARBURST;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARSIZE <= twiddle_rsc_0_4_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARLEN <= twiddle_rsc_0_4_ARLEN;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_ARADDR <= twiddle_rsc_0_4_ARADDR;
  twiddle_rsc_0_4_BRESP <= peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_BRESP;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_WSTRB <= twiddle_rsc_0_4_WSTRB;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_WDATA <= twiddle_rsc_0_4_WDATA;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWREGION <= twiddle_rsc_0_4_AWREGION;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWQOS <= twiddle_rsc_0_4_AWQOS;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWPROT <= twiddle_rsc_0_4_AWPROT;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWCACHE <= twiddle_rsc_0_4_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWBURST <= twiddle_rsc_0_4_AWBURST;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWSIZE <= twiddle_rsc_0_4_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWLEN <= twiddle_rsc_0_4_AWLEN;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_AWADDR <= twiddle_rsc_0_4_AWADDR;
  peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_4_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_4_i_inst_twiddle_rsc_0_4_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_5_i_inst : peaseNTT_core_twiddle_rsc_0_5_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_5_s_tdone => twiddle_rsc_0_5_s_tdone,
      twiddle_rsc_0_5_tr_write_done => twiddle_rsc_0_5_tr_write_done,
      twiddle_rsc_0_5_RREADY => twiddle_rsc_0_5_RREADY,
      twiddle_rsc_0_5_RVALID => twiddle_rsc_0_5_RVALID,
      twiddle_rsc_0_5_RUSER => twiddle_rsc_0_5_RUSER,
      twiddle_rsc_0_5_RLAST => twiddle_rsc_0_5_RLAST,
      twiddle_rsc_0_5_RRESP => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_RRESP,
      twiddle_rsc_0_5_RDATA => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_RDATA,
      twiddle_rsc_0_5_RID => twiddle_rsc_0_5_RID,
      twiddle_rsc_0_5_ARREADY => twiddle_rsc_0_5_ARREADY,
      twiddle_rsc_0_5_ARVALID => twiddle_rsc_0_5_ARVALID,
      twiddle_rsc_0_5_ARUSER => twiddle_rsc_0_5_ARUSER,
      twiddle_rsc_0_5_ARREGION => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARREGION,
      twiddle_rsc_0_5_ARQOS => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARQOS,
      twiddle_rsc_0_5_ARPROT => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARPROT,
      twiddle_rsc_0_5_ARCACHE => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARCACHE,
      twiddle_rsc_0_5_ARLOCK => twiddle_rsc_0_5_ARLOCK,
      twiddle_rsc_0_5_ARBURST => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARBURST,
      twiddle_rsc_0_5_ARSIZE => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARSIZE,
      twiddle_rsc_0_5_ARLEN => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARLEN,
      twiddle_rsc_0_5_ARADDR => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARADDR,
      twiddle_rsc_0_5_ARID => twiddle_rsc_0_5_ARID,
      twiddle_rsc_0_5_BREADY => twiddle_rsc_0_5_BREADY,
      twiddle_rsc_0_5_BVALID => twiddle_rsc_0_5_BVALID,
      twiddle_rsc_0_5_BUSER => twiddle_rsc_0_5_BUSER,
      twiddle_rsc_0_5_BRESP => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_BRESP,
      twiddle_rsc_0_5_BID => twiddle_rsc_0_5_BID,
      twiddle_rsc_0_5_WREADY => twiddle_rsc_0_5_WREADY,
      twiddle_rsc_0_5_WVALID => twiddle_rsc_0_5_WVALID,
      twiddle_rsc_0_5_WUSER => twiddle_rsc_0_5_WUSER,
      twiddle_rsc_0_5_WLAST => twiddle_rsc_0_5_WLAST,
      twiddle_rsc_0_5_WSTRB => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_WSTRB,
      twiddle_rsc_0_5_WDATA => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_WDATA,
      twiddle_rsc_0_5_AWREADY => twiddle_rsc_0_5_AWREADY,
      twiddle_rsc_0_5_AWVALID => twiddle_rsc_0_5_AWVALID,
      twiddle_rsc_0_5_AWUSER => twiddle_rsc_0_5_AWUSER,
      twiddle_rsc_0_5_AWREGION => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWREGION,
      twiddle_rsc_0_5_AWQOS => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWQOS,
      twiddle_rsc_0_5_AWPROT => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWPROT,
      twiddle_rsc_0_5_AWCACHE => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWCACHE,
      twiddle_rsc_0_5_AWLOCK => twiddle_rsc_0_5_AWLOCK,
      twiddle_rsc_0_5_AWBURST => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWBURST,
      twiddle_rsc_0_5_AWSIZE => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWSIZE,
      twiddle_rsc_0_5_AWLEN => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWLEN,
      twiddle_rsc_0_5_AWADDR => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWADDR,
      twiddle_rsc_0_5_AWID => twiddle_rsc_0_5_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_5_i_oswt => reg_twiddle_rsc_0_5_i_oswt_cse,
      twiddle_rsc_0_5_i_wen_comp => twiddle_rsc_0_5_i_wen_comp,
      twiddle_rsc_0_5_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_i_s_raddr_core,
      twiddle_rsc_0_5_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_i_s_din_mxwt
    );
  twiddle_rsc_0_5_RRESP <= peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_RRESP;
  twiddle_rsc_0_5_RDATA <= peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_RDATA;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARREGION <= twiddle_rsc_0_5_ARREGION;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARQOS <= twiddle_rsc_0_5_ARQOS;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARPROT <= twiddle_rsc_0_5_ARPROT;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARCACHE <= twiddle_rsc_0_5_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARBURST <= twiddle_rsc_0_5_ARBURST;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARSIZE <= twiddle_rsc_0_5_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARLEN <= twiddle_rsc_0_5_ARLEN;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_ARADDR <= twiddle_rsc_0_5_ARADDR;
  twiddle_rsc_0_5_BRESP <= peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_BRESP;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_WSTRB <= twiddle_rsc_0_5_WSTRB;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_WDATA <= twiddle_rsc_0_5_WDATA;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWREGION <= twiddle_rsc_0_5_AWREGION;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWQOS <= twiddle_rsc_0_5_AWQOS;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWPROT <= twiddle_rsc_0_5_AWPROT;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWCACHE <= twiddle_rsc_0_5_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWBURST <= twiddle_rsc_0_5_AWBURST;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWSIZE <= twiddle_rsc_0_5_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWLEN <= twiddle_rsc_0_5_AWLEN;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_AWADDR <= twiddle_rsc_0_5_AWADDR;
  peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_5_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_5_i_inst_twiddle_rsc_0_5_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_6_i_inst : peaseNTT_core_twiddle_rsc_0_6_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_6_s_tdone => twiddle_rsc_0_6_s_tdone,
      twiddle_rsc_0_6_tr_write_done => twiddle_rsc_0_6_tr_write_done,
      twiddle_rsc_0_6_RREADY => twiddle_rsc_0_6_RREADY,
      twiddle_rsc_0_6_RVALID => twiddle_rsc_0_6_RVALID,
      twiddle_rsc_0_6_RUSER => twiddle_rsc_0_6_RUSER,
      twiddle_rsc_0_6_RLAST => twiddle_rsc_0_6_RLAST,
      twiddle_rsc_0_6_RRESP => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_RRESP,
      twiddle_rsc_0_6_RDATA => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_RDATA,
      twiddle_rsc_0_6_RID => twiddle_rsc_0_6_RID,
      twiddle_rsc_0_6_ARREADY => twiddle_rsc_0_6_ARREADY,
      twiddle_rsc_0_6_ARVALID => twiddle_rsc_0_6_ARVALID,
      twiddle_rsc_0_6_ARUSER => twiddle_rsc_0_6_ARUSER,
      twiddle_rsc_0_6_ARREGION => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARREGION,
      twiddle_rsc_0_6_ARQOS => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARQOS,
      twiddle_rsc_0_6_ARPROT => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARPROT,
      twiddle_rsc_0_6_ARCACHE => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARCACHE,
      twiddle_rsc_0_6_ARLOCK => twiddle_rsc_0_6_ARLOCK,
      twiddle_rsc_0_6_ARBURST => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARBURST,
      twiddle_rsc_0_6_ARSIZE => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARSIZE,
      twiddle_rsc_0_6_ARLEN => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARLEN,
      twiddle_rsc_0_6_ARADDR => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARADDR,
      twiddle_rsc_0_6_ARID => twiddle_rsc_0_6_ARID,
      twiddle_rsc_0_6_BREADY => twiddle_rsc_0_6_BREADY,
      twiddle_rsc_0_6_BVALID => twiddle_rsc_0_6_BVALID,
      twiddle_rsc_0_6_BUSER => twiddle_rsc_0_6_BUSER,
      twiddle_rsc_0_6_BRESP => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_BRESP,
      twiddle_rsc_0_6_BID => twiddle_rsc_0_6_BID,
      twiddle_rsc_0_6_WREADY => twiddle_rsc_0_6_WREADY,
      twiddle_rsc_0_6_WVALID => twiddle_rsc_0_6_WVALID,
      twiddle_rsc_0_6_WUSER => twiddle_rsc_0_6_WUSER,
      twiddle_rsc_0_6_WLAST => twiddle_rsc_0_6_WLAST,
      twiddle_rsc_0_6_WSTRB => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_WSTRB,
      twiddle_rsc_0_6_WDATA => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_WDATA,
      twiddle_rsc_0_6_AWREADY => twiddle_rsc_0_6_AWREADY,
      twiddle_rsc_0_6_AWVALID => twiddle_rsc_0_6_AWVALID,
      twiddle_rsc_0_6_AWUSER => twiddle_rsc_0_6_AWUSER,
      twiddle_rsc_0_6_AWREGION => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWREGION,
      twiddle_rsc_0_6_AWQOS => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWQOS,
      twiddle_rsc_0_6_AWPROT => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWPROT,
      twiddle_rsc_0_6_AWCACHE => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWCACHE,
      twiddle_rsc_0_6_AWLOCK => twiddle_rsc_0_6_AWLOCK,
      twiddle_rsc_0_6_AWBURST => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWBURST,
      twiddle_rsc_0_6_AWSIZE => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWSIZE,
      twiddle_rsc_0_6_AWLEN => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWLEN,
      twiddle_rsc_0_6_AWADDR => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWADDR,
      twiddle_rsc_0_6_AWID => twiddle_rsc_0_6_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_6_i_oswt => reg_twiddle_rsc_0_6_i_oswt_cse,
      twiddle_rsc_0_6_i_wen_comp => twiddle_rsc_0_6_i_wen_comp,
      twiddle_rsc_0_6_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_i_s_raddr_core,
      twiddle_rsc_0_6_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_i_s_din_mxwt
    );
  twiddle_rsc_0_6_RRESP <= peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_RRESP;
  twiddle_rsc_0_6_RDATA <= peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_RDATA;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARREGION <= twiddle_rsc_0_6_ARREGION;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARQOS <= twiddle_rsc_0_6_ARQOS;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARPROT <= twiddle_rsc_0_6_ARPROT;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARCACHE <= twiddle_rsc_0_6_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARBURST <= twiddle_rsc_0_6_ARBURST;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARSIZE <= twiddle_rsc_0_6_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARLEN <= twiddle_rsc_0_6_ARLEN;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_ARADDR <= twiddle_rsc_0_6_ARADDR;
  twiddle_rsc_0_6_BRESP <= peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_BRESP;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_WSTRB <= twiddle_rsc_0_6_WSTRB;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_WDATA <= twiddle_rsc_0_6_WDATA;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWREGION <= twiddle_rsc_0_6_AWREGION;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWQOS <= twiddle_rsc_0_6_AWQOS;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWPROT <= twiddle_rsc_0_6_AWPROT;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWCACHE <= twiddle_rsc_0_6_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWBURST <= twiddle_rsc_0_6_AWBURST;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWSIZE <= twiddle_rsc_0_6_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWLEN <= twiddle_rsc_0_6_AWLEN;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_AWADDR <= twiddle_rsc_0_6_AWADDR;
  peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_6_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_6_i_inst_twiddle_rsc_0_6_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_7_i_inst : peaseNTT_core_twiddle_rsc_0_7_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_7_s_tdone => twiddle_rsc_0_7_s_tdone,
      twiddle_rsc_0_7_tr_write_done => twiddle_rsc_0_7_tr_write_done,
      twiddle_rsc_0_7_RREADY => twiddle_rsc_0_7_RREADY,
      twiddle_rsc_0_7_RVALID => twiddle_rsc_0_7_RVALID,
      twiddle_rsc_0_7_RUSER => twiddle_rsc_0_7_RUSER,
      twiddle_rsc_0_7_RLAST => twiddle_rsc_0_7_RLAST,
      twiddle_rsc_0_7_RRESP => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_RRESP,
      twiddle_rsc_0_7_RDATA => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_RDATA,
      twiddle_rsc_0_7_RID => twiddle_rsc_0_7_RID,
      twiddle_rsc_0_7_ARREADY => twiddle_rsc_0_7_ARREADY,
      twiddle_rsc_0_7_ARVALID => twiddle_rsc_0_7_ARVALID,
      twiddle_rsc_0_7_ARUSER => twiddle_rsc_0_7_ARUSER,
      twiddle_rsc_0_7_ARREGION => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARREGION,
      twiddle_rsc_0_7_ARQOS => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARQOS,
      twiddle_rsc_0_7_ARPROT => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARPROT,
      twiddle_rsc_0_7_ARCACHE => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARCACHE,
      twiddle_rsc_0_7_ARLOCK => twiddle_rsc_0_7_ARLOCK,
      twiddle_rsc_0_7_ARBURST => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARBURST,
      twiddle_rsc_0_7_ARSIZE => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARSIZE,
      twiddle_rsc_0_7_ARLEN => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARLEN,
      twiddle_rsc_0_7_ARADDR => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARADDR,
      twiddle_rsc_0_7_ARID => twiddle_rsc_0_7_ARID,
      twiddle_rsc_0_7_BREADY => twiddle_rsc_0_7_BREADY,
      twiddle_rsc_0_7_BVALID => twiddle_rsc_0_7_BVALID,
      twiddle_rsc_0_7_BUSER => twiddle_rsc_0_7_BUSER,
      twiddle_rsc_0_7_BRESP => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_BRESP,
      twiddle_rsc_0_7_BID => twiddle_rsc_0_7_BID,
      twiddle_rsc_0_7_WREADY => twiddle_rsc_0_7_WREADY,
      twiddle_rsc_0_7_WVALID => twiddle_rsc_0_7_WVALID,
      twiddle_rsc_0_7_WUSER => twiddle_rsc_0_7_WUSER,
      twiddle_rsc_0_7_WLAST => twiddle_rsc_0_7_WLAST,
      twiddle_rsc_0_7_WSTRB => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_WSTRB,
      twiddle_rsc_0_7_WDATA => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_WDATA,
      twiddle_rsc_0_7_AWREADY => twiddle_rsc_0_7_AWREADY,
      twiddle_rsc_0_7_AWVALID => twiddle_rsc_0_7_AWVALID,
      twiddle_rsc_0_7_AWUSER => twiddle_rsc_0_7_AWUSER,
      twiddle_rsc_0_7_AWREGION => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWREGION,
      twiddle_rsc_0_7_AWQOS => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWQOS,
      twiddle_rsc_0_7_AWPROT => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWPROT,
      twiddle_rsc_0_7_AWCACHE => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWCACHE,
      twiddle_rsc_0_7_AWLOCK => twiddle_rsc_0_7_AWLOCK,
      twiddle_rsc_0_7_AWBURST => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWBURST,
      twiddle_rsc_0_7_AWSIZE => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWSIZE,
      twiddle_rsc_0_7_AWLEN => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWLEN,
      twiddle_rsc_0_7_AWADDR => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWADDR,
      twiddle_rsc_0_7_AWID => twiddle_rsc_0_7_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_7_i_oswt => reg_twiddle_rsc_0_7_i_oswt_cse,
      twiddle_rsc_0_7_i_wen_comp => twiddle_rsc_0_7_i_wen_comp,
      twiddle_rsc_0_7_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_i_s_raddr_core,
      twiddle_rsc_0_7_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_i_s_din_mxwt
    );
  twiddle_rsc_0_7_RRESP <= peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_RRESP;
  twiddle_rsc_0_7_RDATA <= peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_RDATA;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARREGION <= twiddle_rsc_0_7_ARREGION;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARQOS <= twiddle_rsc_0_7_ARQOS;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARPROT <= twiddle_rsc_0_7_ARPROT;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARCACHE <= twiddle_rsc_0_7_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARBURST <= twiddle_rsc_0_7_ARBURST;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARSIZE <= twiddle_rsc_0_7_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARLEN <= twiddle_rsc_0_7_ARLEN;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_ARADDR <= twiddle_rsc_0_7_ARADDR;
  twiddle_rsc_0_7_BRESP <= peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_BRESP;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_WSTRB <= twiddle_rsc_0_7_WSTRB;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_WDATA <= twiddle_rsc_0_7_WDATA;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWREGION <= twiddle_rsc_0_7_AWREGION;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWQOS <= twiddle_rsc_0_7_AWQOS;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWPROT <= twiddle_rsc_0_7_AWPROT;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWCACHE <= twiddle_rsc_0_7_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWBURST <= twiddle_rsc_0_7_AWBURST;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWSIZE <= twiddle_rsc_0_7_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWLEN <= twiddle_rsc_0_7_AWLEN;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_AWADDR <= twiddle_rsc_0_7_AWADDR;
  peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_7_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_7_i_inst_twiddle_rsc_0_7_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_8_i_inst : peaseNTT_core_twiddle_rsc_0_8_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_8_s_tdone => twiddle_rsc_0_8_s_tdone,
      twiddle_rsc_0_8_tr_write_done => twiddle_rsc_0_8_tr_write_done,
      twiddle_rsc_0_8_RREADY => twiddle_rsc_0_8_RREADY,
      twiddle_rsc_0_8_RVALID => twiddle_rsc_0_8_RVALID,
      twiddle_rsc_0_8_RUSER => twiddle_rsc_0_8_RUSER,
      twiddle_rsc_0_8_RLAST => twiddle_rsc_0_8_RLAST,
      twiddle_rsc_0_8_RRESP => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_RRESP,
      twiddle_rsc_0_8_RDATA => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_RDATA,
      twiddle_rsc_0_8_RID => twiddle_rsc_0_8_RID,
      twiddle_rsc_0_8_ARREADY => twiddle_rsc_0_8_ARREADY,
      twiddle_rsc_0_8_ARVALID => twiddle_rsc_0_8_ARVALID,
      twiddle_rsc_0_8_ARUSER => twiddle_rsc_0_8_ARUSER,
      twiddle_rsc_0_8_ARREGION => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARREGION,
      twiddle_rsc_0_8_ARQOS => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARQOS,
      twiddle_rsc_0_8_ARPROT => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARPROT,
      twiddle_rsc_0_8_ARCACHE => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARCACHE,
      twiddle_rsc_0_8_ARLOCK => twiddle_rsc_0_8_ARLOCK,
      twiddle_rsc_0_8_ARBURST => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARBURST,
      twiddle_rsc_0_8_ARSIZE => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARSIZE,
      twiddle_rsc_0_8_ARLEN => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARLEN,
      twiddle_rsc_0_8_ARADDR => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARADDR,
      twiddle_rsc_0_8_ARID => twiddle_rsc_0_8_ARID,
      twiddle_rsc_0_8_BREADY => twiddle_rsc_0_8_BREADY,
      twiddle_rsc_0_8_BVALID => twiddle_rsc_0_8_BVALID,
      twiddle_rsc_0_8_BUSER => twiddle_rsc_0_8_BUSER,
      twiddle_rsc_0_8_BRESP => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_BRESP,
      twiddle_rsc_0_8_BID => twiddle_rsc_0_8_BID,
      twiddle_rsc_0_8_WREADY => twiddle_rsc_0_8_WREADY,
      twiddle_rsc_0_8_WVALID => twiddle_rsc_0_8_WVALID,
      twiddle_rsc_0_8_WUSER => twiddle_rsc_0_8_WUSER,
      twiddle_rsc_0_8_WLAST => twiddle_rsc_0_8_WLAST,
      twiddle_rsc_0_8_WSTRB => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_WSTRB,
      twiddle_rsc_0_8_WDATA => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_WDATA,
      twiddle_rsc_0_8_AWREADY => twiddle_rsc_0_8_AWREADY,
      twiddle_rsc_0_8_AWVALID => twiddle_rsc_0_8_AWVALID,
      twiddle_rsc_0_8_AWUSER => twiddle_rsc_0_8_AWUSER,
      twiddle_rsc_0_8_AWREGION => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWREGION,
      twiddle_rsc_0_8_AWQOS => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWQOS,
      twiddle_rsc_0_8_AWPROT => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWPROT,
      twiddle_rsc_0_8_AWCACHE => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWCACHE,
      twiddle_rsc_0_8_AWLOCK => twiddle_rsc_0_8_AWLOCK,
      twiddle_rsc_0_8_AWBURST => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWBURST,
      twiddle_rsc_0_8_AWSIZE => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWSIZE,
      twiddle_rsc_0_8_AWLEN => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWLEN,
      twiddle_rsc_0_8_AWADDR => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWADDR,
      twiddle_rsc_0_8_AWID => twiddle_rsc_0_8_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_8_i_oswt => reg_twiddle_rsc_0_8_i_oswt_cse,
      twiddle_rsc_0_8_i_wen_comp => twiddle_rsc_0_8_i_wen_comp,
      twiddle_rsc_0_8_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_i_s_raddr_core,
      twiddle_rsc_0_8_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_i_s_din_mxwt
    );
  twiddle_rsc_0_8_RRESP <= peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_RRESP;
  twiddle_rsc_0_8_RDATA <= peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_RDATA;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARREGION <= twiddle_rsc_0_8_ARREGION;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARQOS <= twiddle_rsc_0_8_ARQOS;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARPROT <= twiddle_rsc_0_8_ARPROT;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARCACHE <= twiddle_rsc_0_8_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARBURST <= twiddle_rsc_0_8_ARBURST;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARSIZE <= twiddle_rsc_0_8_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARLEN <= twiddle_rsc_0_8_ARLEN;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_ARADDR <= twiddle_rsc_0_8_ARADDR;
  twiddle_rsc_0_8_BRESP <= peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_BRESP;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_WSTRB <= twiddle_rsc_0_8_WSTRB;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_WDATA <= twiddle_rsc_0_8_WDATA;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWREGION <= twiddle_rsc_0_8_AWREGION;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWQOS <= twiddle_rsc_0_8_AWQOS;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWPROT <= twiddle_rsc_0_8_AWPROT;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWCACHE <= twiddle_rsc_0_8_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWBURST <= twiddle_rsc_0_8_AWBURST;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWSIZE <= twiddle_rsc_0_8_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWLEN <= twiddle_rsc_0_8_AWLEN;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_AWADDR <= twiddle_rsc_0_8_AWADDR;
  peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_8_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_8_i_inst_twiddle_rsc_0_8_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_9_i_inst : peaseNTT_core_twiddle_rsc_0_9_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_9_s_tdone => twiddle_rsc_0_9_s_tdone,
      twiddle_rsc_0_9_tr_write_done => twiddle_rsc_0_9_tr_write_done,
      twiddle_rsc_0_9_RREADY => twiddle_rsc_0_9_RREADY,
      twiddle_rsc_0_9_RVALID => twiddle_rsc_0_9_RVALID,
      twiddle_rsc_0_9_RUSER => twiddle_rsc_0_9_RUSER,
      twiddle_rsc_0_9_RLAST => twiddle_rsc_0_9_RLAST,
      twiddle_rsc_0_9_RRESP => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_RRESP,
      twiddle_rsc_0_9_RDATA => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_RDATA,
      twiddle_rsc_0_9_RID => twiddle_rsc_0_9_RID,
      twiddle_rsc_0_9_ARREADY => twiddle_rsc_0_9_ARREADY,
      twiddle_rsc_0_9_ARVALID => twiddle_rsc_0_9_ARVALID,
      twiddle_rsc_0_9_ARUSER => twiddle_rsc_0_9_ARUSER,
      twiddle_rsc_0_9_ARREGION => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARREGION,
      twiddle_rsc_0_9_ARQOS => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARQOS,
      twiddle_rsc_0_9_ARPROT => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARPROT,
      twiddle_rsc_0_9_ARCACHE => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARCACHE,
      twiddle_rsc_0_9_ARLOCK => twiddle_rsc_0_9_ARLOCK,
      twiddle_rsc_0_9_ARBURST => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARBURST,
      twiddle_rsc_0_9_ARSIZE => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARSIZE,
      twiddle_rsc_0_9_ARLEN => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARLEN,
      twiddle_rsc_0_9_ARADDR => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARADDR,
      twiddle_rsc_0_9_ARID => twiddle_rsc_0_9_ARID,
      twiddle_rsc_0_9_BREADY => twiddle_rsc_0_9_BREADY,
      twiddle_rsc_0_9_BVALID => twiddle_rsc_0_9_BVALID,
      twiddle_rsc_0_9_BUSER => twiddle_rsc_0_9_BUSER,
      twiddle_rsc_0_9_BRESP => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_BRESP,
      twiddle_rsc_0_9_BID => twiddle_rsc_0_9_BID,
      twiddle_rsc_0_9_WREADY => twiddle_rsc_0_9_WREADY,
      twiddle_rsc_0_9_WVALID => twiddle_rsc_0_9_WVALID,
      twiddle_rsc_0_9_WUSER => twiddle_rsc_0_9_WUSER,
      twiddle_rsc_0_9_WLAST => twiddle_rsc_0_9_WLAST,
      twiddle_rsc_0_9_WSTRB => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_WSTRB,
      twiddle_rsc_0_9_WDATA => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_WDATA,
      twiddle_rsc_0_9_AWREADY => twiddle_rsc_0_9_AWREADY,
      twiddle_rsc_0_9_AWVALID => twiddle_rsc_0_9_AWVALID,
      twiddle_rsc_0_9_AWUSER => twiddle_rsc_0_9_AWUSER,
      twiddle_rsc_0_9_AWREGION => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWREGION,
      twiddle_rsc_0_9_AWQOS => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWQOS,
      twiddle_rsc_0_9_AWPROT => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWPROT,
      twiddle_rsc_0_9_AWCACHE => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWCACHE,
      twiddle_rsc_0_9_AWLOCK => twiddle_rsc_0_9_AWLOCK,
      twiddle_rsc_0_9_AWBURST => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWBURST,
      twiddle_rsc_0_9_AWSIZE => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWSIZE,
      twiddle_rsc_0_9_AWLEN => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWLEN,
      twiddle_rsc_0_9_AWADDR => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWADDR,
      twiddle_rsc_0_9_AWID => twiddle_rsc_0_9_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_9_i_oswt => reg_twiddle_rsc_0_1_i_oswt_cse,
      twiddle_rsc_0_9_i_wen_comp => twiddle_rsc_0_9_i_wen_comp,
      twiddle_rsc_0_9_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_i_s_raddr_core,
      twiddle_rsc_0_9_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_i_s_din_mxwt
    );
  twiddle_rsc_0_9_RRESP <= peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_RRESP;
  twiddle_rsc_0_9_RDATA <= peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_RDATA;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARREGION <= twiddle_rsc_0_9_ARREGION;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARQOS <= twiddle_rsc_0_9_ARQOS;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARPROT <= twiddle_rsc_0_9_ARPROT;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARCACHE <= twiddle_rsc_0_9_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARBURST <= twiddle_rsc_0_9_ARBURST;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARSIZE <= twiddle_rsc_0_9_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARLEN <= twiddle_rsc_0_9_ARLEN;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_ARADDR <= twiddle_rsc_0_9_ARADDR;
  twiddle_rsc_0_9_BRESP <= peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_BRESP;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_WSTRB <= twiddle_rsc_0_9_WSTRB;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_WDATA <= twiddle_rsc_0_9_WDATA;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWREGION <= twiddle_rsc_0_9_AWREGION;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWQOS <= twiddle_rsc_0_9_AWQOS;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWPROT <= twiddle_rsc_0_9_AWPROT;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWCACHE <= twiddle_rsc_0_9_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWBURST <= twiddle_rsc_0_9_AWBURST;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWSIZE <= twiddle_rsc_0_9_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWLEN <= twiddle_rsc_0_9_AWLEN;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_AWADDR <= twiddle_rsc_0_9_AWADDR;
  peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_9_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_9_i_inst_twiddle_rsc_0_9_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_10_i_inst : peaseNTT_core_twiddle_rsc_0_10_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_10_s_tdone => twiddle_rsc_0_10_s_tdone,
      twiddle_rsc_0_10_tr_write_done => twiddle_rsc_0_10_tr_write_done,
      twiddle_rsc_0_10_RREADY => twiddle_rsc_0_10_RREADY,
      twiddle_rsc_0_10_RVALID => twiddle_rsc_0_10_RVALID,
      twiddle_rsc_0_10_RUSER => twiddle_rsc_0_10_RUSER,
      twiddle_rsc_0_10_RLAST => twiddle_rsc_0_10_RLAST,
      twiddle_rsc_0_10_RRESP => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_RRESP,
      twiddle_rsc_0_10_RDATA => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_RDATA,
      twiddle_rsc_0_10_RID => twiddle_rsc_0_10_RID,
      twiddle_rsc_0_10_ARREADY => twiddle_rsc_0_10_ARREADY,
      twiddle_rsc_0_10_ARVALID => twiddle_rsc_0_10_ARVALID,
      twiddle_rsc_0_10_ARUSER => twiddle_rsc_0_10_ARUSER,
      twiddle_rsc_0_10_ARREGION => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARREGION,
      twiddle_rsc_0_10_ARQOS => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARQOS,
      twiddle_rsc_0_10_ARPROT => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARPROT,
      twiddle_rsc_0_10_ARCACHE => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARCACHE,
      twiddle_rsc_0_10_ARLOCK => twiddle_rsc_0_10_ARLOCK,
      twiddle_rsc_0_10_ARBURST => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARBURST,
      twiddle_rsc_0_10_ARSIZE => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARSIZE,
      twiddle_rsc_0_10_ARLEN => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARLEN,
      twiddle_rsc_0_10_ARADDR => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARADDR,
      twiddle_rsc_0_10_ARID => twiddle_rsc_0_10_ARID,
      twiddle_rsc_0_10_BREADY => twiddle_rsc_0_10_BREADY,
      twiddle_rsc_0_10_BVALID => twiddle_rsc_0_10_BVALID,
      twiddle_rsc_0_10_BUSER => twiddle_rsc_0_10_BUSER,
      twiddle_rsc_0_10_BRESP => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_BRESP,
      twiddle_rsc_0_10_BID => twiddle_rsc_0_10_BID,
      twiddle_rsc_0_10_WREADY => twiddle_rsc_0_10_WREADY,
      twiddle_rsc_0_10_WVALID => twiddle_rsc_0_10_WVALID,
      twiddle_rsc_0_10_WUSER => twiddle_rsc_0_10_WUSER,
      twiddle_rsc_0_10_WLAST => twiddle_rsc_0_10_WLAST,
      twiddle_rsc_0_10_WSTRB => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_WSTRB,
      twiddle_rsc_0_10_WDATA => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_WDATA,
      twiddle_rsc_0_10_AWREADY => twiddle_rsc_0_10_AWREADY,
      twiddle_rsc_0_10_AWVALID => twiddle_rsc_0_10_AWVALID,
      twiddle_rsc_0_10_AWUSER => twiddle_rsc_0_10_AWUSER,
      twiddle_rsc_0_10_AWREGION => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWREGION,
      twiddle_rsc_0_10_AWQOS => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWQOS,
      twiddle_rsc_0_10_AWPROT => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWPROT,
      twiddle_rsc_0_10_AWCACHE => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWCACHE,
      twiddle_rsc_0_10_AWLOCK => twiddle_rsc_0_10_AWLOCK,
      twiddle_rsc_0_10_AWBURST => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWBURST,
      twiddle_rsc_0_10_AWSIZE => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWSIZE,
      twiddle_rsc_0_10_AWLEN => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWLEN,
      twiddle_rsc_0_10_AWADDR => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWADDR,
      twiddle_rsc_0_10_AWID => twiddle_rsc_0_10_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_10_i_oswt => reg_twiddle_rsc_0_2_i_oswt_cse,
      twiddle_rsc_0_10_i_wen_comp => twiddle_rsc_0_10_i_wen_comp,
      twiddle_rsc_0_10_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_i_s_raddr_core,
      twiddle_rsc_0_10_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_i_s_din_mxwt
    );
  twiddle_rsc_0_10_RRESP <= peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_RRESP;
  twiddle_rsc_0_10_RDATA <= peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_RDATA;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARREGION <= twiddle_rsc_0_10_ARREGION;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARQOS <= twiddle_rsc_0_10_ARQOS;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARPROT <= twiddle_rsc_0_10_ARPROT;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARCACHE <= twiddle_rsc_0_10_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARBURST <= twiddle_rsc_0_10_ARBURST;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARSIZE <= twiddle_rsc_0_10_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARLEN <= twiddle_rsc_0_10_ARLEN;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_ARADDR <= twiddle_rsc_0_10_ARADDR;
  twiddle_rsc_0_10_BRESP <= peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_BRESP;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_WSTRB <= twiddle_rsc_0_10_WSTRB;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_WDATA <= twiddle_rsc_0_10_WDATA;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWREGION <= twiddle_rsc_0_10_AWREGION;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWQOS <= twiddle_rsc_0_10_AWQOS;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWPROT <= twiddle_rsc_0_10_AWPROT;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWCACHE <= twiddle_rsc_0_10_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWBURST <= twiddle_rsc_0_10_AWBURST;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWSIZE <= twiddle_rsc_0_10_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWLEN <= twiddle_rsc_0_10_AWLEN;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_AWADDR <= twiddle_rsc_0_10_AWADDR;
  peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_10_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_10_i_inst_twiddle_rsc_0_10_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_11_i_inst : peaseNTT_core_twiddle_rsc_0_11_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_11_s_tdone => twiddle_rsc_0_11_s_tdone,
      twiddle_rsc_0_11_tr_write_done => twiddle_rsc_0_11_tr_write_done,
      twiddle_rsc_0_11_RREADY => twiddle_rsc_0_11_RREADY,
      twiddle_rsc_0_11_RVALID => twiddle_rsc_0_11_RVALID,
      twiddle_rsc_0_11_RUSER => twiddle_rsc_0_11_RUSER,
      twiddle_rsc_0_11_RLAST => twiddle_rsc_0_11_RLAST,
      twiddle_rsc_0_11_RRESP => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_RRESP,
      twiddle_rsc_0_11_RDATA => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_RDATA,
      twiddle_rsc_0_11_RID => twiddle_rsc_0_11_RID,
      twiddle_rsc_0_11_ARREADY => twiddle_rsc_0_11_ARREADY,
      twiddle_rsc_0_11_ARVALID => twiddle_rsc_0_11_ARVALID,
      twiddle_rsc_0_11_ARUSER => twiddle_rsc_0_11_ARUSER,
      twiddle_rsc_0_11_ARREGION => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARREGION,
      twiddle_rsc_0_11_ARQOS => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARQOS,
      twiddle_rsc_0_11_ARPROT => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARPROT,
      twiddle_rsc_0_11_ARCACHE => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARCACHE,
      twiddle_rsc_0_11_ARLOCK => twiddle_rsc_0_11_ARLOCK,
      twiddle_rsc_0_11_ARBURST => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARBURST,
      twiddle_rsc_0_11_ARSIZE => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARSIZE,
      twiddle_rsc_0_11_ARLEN => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARLEN,
      twiddle_rsc_0_11_ARADDR => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARADDR,
      twiddle_rsc_0_11_ARID => twiddle_rsc_0_11_ARID,
      twiddle_rsc_0_11_BREADY => twiddle_rsc_0_11_BREADY,
      twiddle_rsc_0_11_BVALID => twiddle_rsc_0_11_BVALID,
      twiddle_rsc_0_11_BUSER => twiddle_rsc_0_11_BUSER,
      twiddle_rsc_0_11_BRESP => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_BRESP,
      twiddle_rsc_0_11_BID => twiddle_rsc_0_11_BID,
      twiddle_rsc_0_11_WREADY => twiddle_rsc_0_11_WREADY,
      twiddle_rsc_0_11_WVALID => twiddle_rsc_0_11_WVALID,
      twiddle_rsc_0_11_WUSER => twiddle_rsc_0_11_WUSER,
      twiddle_rsc_0_11_WLAST => twiddle_rsc_0_11_WLAST,
      twiddle_rsc_0_11_WSTRB => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_WSTRB,
      twiddle_rsc_0_11_WDATA => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_WDATA,
      twiddle_rsc_0_11_AWREADY => twiddle_rsc_0_11_AWREADY,
      twiddle_rsc_0_11_AWVALID => twiddle_rsc_0_11_AWVALID,
      twiddle_rsc_0_11_AWUSER => twiddle_rsc_0_11_AWUSER,
      twiddle_rsc_0_11_AWREGION => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWREGION,
      twiddle_rsc_0_11_AWQOS => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWQOS,
      twiddle_rsc_0_11_AWPROT => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWPROT,
      twiddle_rsc_0_11_AWCACHE => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWCACHE,
      twiddle_rsc_0_11_AWLOCK => twiddle_rsc_0_11_AWLOCK,
      twiddle_rsc_0_11_AWBURST => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWBURST,
      twiddle_rsc_0_11_AWSIZE => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWSIZE,
      twiddle_rsc_0_11_AWLEN => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWLEN,
      twiddle_rsc_0_11_AWADDR => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWADDR,
      twiddle_rsc_0_11_AWID => twiddle_rsc_0_11_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_11_i_oswt => reg_twiddle_rsc_0_3_i_oswt_cse,
      twiddle_rsc_0_11_i_wen_comp => twiddle_rsc_0_11_i_wen_comp,
      twiddle_rsc_0_11_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_i_s_raddr_core,
      twiddle_rsc_0_11_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_i_s_din_mxwt
    );
  twiddle_rsc_0_11_RRESP <= peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_RRESP;
  twiddle_rsc_0_11_RDATA <= peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_RDATA;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARREGION <= twiddle_rsc_0_11_ARREGION;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARQOS <= twiddle_rsc_0_11_ARQOS;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARPROT <= twiddle_rsc_0_11_ARPROT;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARCACHE <= twiddle_rsc_0_11_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARBURST <= twiddle_rsc_0_11_ARBURST;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARSIZE <= twiddle_rsc_0_11_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARLEN <= twiddle_rsc_0_11_ARLEN;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_ARADDR <= twiddle_rsc_0_11_ARADDR;
  twiddle_rsc_0_11_BRESP <= peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_BRESP;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_WSTRB <= twiddle_rsc_0_11_WSTRB;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_WDATA <= twiddle_rsc_0_11_WDATA;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWREGION <= twiddle_rsc_0_11_AWREGION;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWQOS <= twiddle_rsc_0_11_AWQOS;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWPROT <= twiddle_rsc_0_11_AWPROT;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWCACHE <= twiddle_rsc_0_11_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWBURST <= twiddle_rsc_0_11_AWBURST;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWSIZE <= twiddle_rsc_0_11_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWLEN <= twiddle_rsc_0_11_AWLEN;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_AWADDR <= twiddle_rsc_0_11_AWADDR;
  peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_11_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_11_i_inst_twiddle_rsc_0_11_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_12_i_inst : peaseNTT_core_twiddle_rsc_0_12_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_12_s_tdone => twiddle_rsc_0_12_s_tdone,
      twiddle_rsc_0_12_tr_write_done => twiddle_rsc_0_12_tr_write_done,
      twiddle_rsc_0_12_RREADY => twiddle_rsc_0_12_RREADY,
      twiddle_rsc_0_12_RVALID => twiddle_rsc_0_12_RVALID,
      twiddle_rsc_0_12_RUSER => twiddle_rsc_0_12_RUSER,
      twiddle_rsc_0_12_RLAST => twiddle_rsc_0_12_RLAST,
      twiddle_rsc_0_12_RRESP => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_RRESP,
      twiddle_rsc_0_12_RDATA => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_RDATA,
      twiddle_rsc_0_12_RID => twiddle_rsc_0_12_RID,
      twiddle_rsc_0_12_ARREADY => twiddle_rsc_0_12_ARREADY,
      twiddle_rsc_0_12_ARVALID => twiddle_rsc_0_12_ARVALID,
      twiddle_rsc_0_12_ARUSER => twiddle_rsc_0_12_ARUSER,
      twiddle_rsc_0_12_ARREGION => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARREGION,
      twiddle_rsc_0_12_ARQOS => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARQOS,
      twiddle_rsc_0_12_ARPROT => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARPROT,
      twiddle_rsc_0_12_ARCACHE => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARCACHE,
      twiddle_rsc_0_12_ARLOCK => twiddle_rsc_0_12_ARLOCK,
      twiddle_rsc_0_12_ARBURST => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARBURST,
      twiddle_rsc_0_12_ARSIZE => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARSIZE,
      twiddle_rsc_0_12_ARLEN => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARLEN,
      twiddle_rsc_0_12_ARADDR => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARADDR,
      twiddle_rsc_0_12_ARID => twiddle_rsc_0_12_ARID,
      twiddle_rsc_0_12_BREADY => twiddle_rsc_0_12_BREADY,
      twiddle_rsc_0_12_BVALID => twiddle_rsc_0_12_BVALID,
      twiddle_rsc_0_12_BUSER => twiddle_rsc_0_12_BUSER,
      twiddle_rsc_0_12_BRESP => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_BRESP,
      twiddle_rsc_0_12_BID => twiddle_rsc_0_12_BID,
      twiddle_rsc_0_12_WREADY => twiddle_rsc_0_12_WREADY,
      twiddle_rsc_0_12_WVALID => twiddle_rsc_0_12_WVALID,
      twiddle_rsc_0_12_WUSER => twiddle_rsc_0_12_WUSER,
      twiddle_rsc_0_12_WLAST => twiddle_rsc_0_12_WLAST,
      twiddle_rsc_0_12_WSTRB => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_WSTRB,
      twiddle_rsc_0_12_WDATA => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_WDATA,
      twiddle_rsc_0_12_AWREADY => twiddle_rsc_0_12_AWREADY,
      twiddle_rsc_0_12_AWVALID => twiddle_rsc_0_12_AWVALID,
      twiddle_rsc_0_12_AWUSER => twiddle_rsc_0_12_AWUSER,
      twiddle_rsc_0_12_AWREGION => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWREGION,
      twiddle_rsc_0_12_AWQOS => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWQOS,
      twiddle_rsc_0_12_AWPROT => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWPROT,
      twiddle_rsc_0_12_AWCACHE => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWCACHE,
      twiddle_rsc_0_12_AWLOCK => twiddle_rsc_0_12_AWLOCK,
      twiddle_rsc_0_12_AWBURST => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWBURST,
      twiddle_rsc_0_12_AWSIZE => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWSIZE,
      twiddle_rsc_0_12_AWLEN => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWLEN,
      twiddle_rsc_0_12_AWADDR => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWADDR,
      twiddle_rsc_0_12_AWID => twiddle_rsc_0_12_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_12_i_oswt => reg_twiddle_rsc_0_4_i_oswt_cse,
      twiddle_rsc_0_12_i_wen_comp => twiddle_rsc_0_12_i_wen_comp,
      twiddle_rsc_0_12_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_i_s_raddr_core,
      twiddle_rsc_0_12_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_i_s_din_mxwt
    );
  twiddle_rsc_0_12_RRESP <= peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_RRESP;
  twiddle_rsc_0_12_RDATA <= peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_RDATA;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARREGION <= twiddle_rsc_0_12_ARREGION;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARQOS <= twiddle_rsc_0_12_ARQOS;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARPROT <= twiddle_rsc_0_12_ARPROT;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARCACHE <= twiddle_rsc_0_12_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARBURST <= twiddle_rsc_0_12_ARBURST;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARSIZE <= twiddle_rsc_0_12_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARLEN <= twiddle_rsc_0_12_ARLEN;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_ARADDR <= twiddle_rsc_0_12_ARADDR;
  twiddle_rsc_0_12_BRESP <= peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_BRESP;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_WSTRB <= twiddle_rsc_0_12_WSTRB;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_WDATA <= twiddle_rsc_0_12_WDATA;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWREGION <= twiddle_rsc_0_12_AWREGION;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWQOS <= twiddle_rsc_0_12_AWQOS;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWPROT <= twiddle_rsc_0_12_AWPROT;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWCACHE <= twiddle_rsc_0_12_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWBURST <= twiddle_rsc_0_12_AWBURST;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWSIZE <= twiddle_rsc_0_12_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWLEN <= twiddle_rsc_0_12_AWLEN;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_AWADDR <= twiddle_rsc_0_12_AWADDR;
  peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_12_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_12_i_inst_twiddle_rsc_0_12_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_13_i_inst : peaseNTT_core_twiddle_rsc_0_13_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_13_s_tdone => twiddle_rsc_0_13_s_tdone,
      twiddle_rsc_0_13_tr_write_done => twiddle_rsc_0_13_tr_write_done,
      twiddle_rsc_0_13_RREADY => twiddle_rsc_0_13_RREADY,
      twiddle_rsc_0_13_RVALID => twiddle_rsc_0_13_RVALID,
      twiddle_rsc_0_13_RUSER => twiddle_rsc_0_13_RUSER,
      twiddle_rsc_0_13_RLAST => twiddle_rsc_0_13_RLAST,
      twiddle_rsc_0_13_RRESP => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_RRESP,
      twiddle_rsc_0_13_RDATA => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_RDATA,
      twiddle_rsc_0_13_RID => twiddle_rsc_0_13_RID,
      twiddle_rsc_0_13_ARREADY => twiddle_rsc_0_13_ARREADY,
      twiddle_rsc_0_13_ARVALID => twiddle_rsc_0_13_ARVALID,
      twiddle_rsc_0_13_ARUSER => twiddle_rsc_0_13_ARUSER,
      twiddle_rsc_0_13_ARREGION => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARREGION,
      twiddle_rsc_0_13_ARQOS => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARQOS,
      twiddle_rsc_0_13_ARPROT => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARPROT,
      twiddle_rsc_0_13_ARCACHE => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARCACHE,
      twiddle_rsc_0_13_ARLOCK => twiddle_rsc_0_13_ARLOCK,
      twiddle_rsc_0_13_ARBURST => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARBURST,
      twiddle_rsc_0_13_ARSIZE => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARSIZE,
      twiddle_rsc_0_13_ARLEN => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARLEN,
      twiddle_rsc_0_13_ARADDR => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARADDR,
      twiddle_rsc_0_13_ARID => twiddle_rsc_0_13_ARID,
      twiddle_rsc_0_13_BREADY => twiddle_rsc_0_13_BREADY,
      twiddle_rsc_0_13_BVALID => twiddle_rsc_0_13_BVALID,
      twiddle_rsc_0_13_BUSER => twiddle_rsc_0_13_BUSER,
      twiddle_rsc_0_13_BRESP => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_BRESP,
      twiddle_rsc_0_13_BID => twiddle_rsc_0_13_BID,
      twiddle_rsc_0_13_WREADY => twiddle_rsc_0_13_WREADY,
      twiddle_rsc_0_13_WVALID => twiddle_rsc_0_13_WVALID,
      twiddle_rsc_0_13_WUSER => twiddle_rsc_0_13_WUSER,
      twiddle_rsc_0_13_WLAST => twiddle_rsc_0_13_WLAST,
      twiddle_rsc_0_13_WSTRB => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_WSTRB,
      twiddle_rsc_0_13_WDATA => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_WDATA,
      twiddle_rsc_0_13_AWREADY => twiddle_rsc_0_13_AWREADY,
      twiddle_rsc_0_13_AWVALID => twiddle_rsc_0_13_AWVALID,
      twiddle_rsc_0_13_AWUSER => twiddle_rsc_0_13_AWUSER,
      twiddle_rsc_0_13_AWREGION => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWREGION,
      twiddle_rsc_0_13_AWQOS => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWQOS,
      twiddle_rsc_0_13_AWPROT => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWPROT,
      twiddle_rsc_0_13_AWCACHE => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWCACHE,
      twiddle_rsc_0_13_AWLOCK => twiddle_rsc_0_13_AWLOCK,
      twiddle_rsc_0_13_AWBURST => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWBURST,
      twiddle_rsc_0_13_AWSIZE => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWSIZE,
      twiddle_rsc_0_13_AWLEN => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWLEN,
      twiddle_rsc_0_13_AWADDR => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWADDR,
      twiddle_rsc_0_13_AWID => twiddle_rsc_0_13_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_13_i_oswt => reg_twiddle_rsc_0_5_i_oswt_cse,
      twiddle_rsc_0_13_i_wen_comp => twiddle_rsc_0_13_i_wen_comp,
      twiddle_rsc_0_13_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_i_s_raddr_core,
      twiddle_rsc_0_13_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_i_s_din_mxwt
    );
  twiddle_rsc_0_13_RRESP <= peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_RRESP;
  twiddle_rsc_0_13_RDATA <= peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_RDATA;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARREGION <= twiddle_rsc_0_13_ARREGION;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARQOS <= twiddle_rsc_0_13_ARQOS;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARPROT <= twiddle_rsc_0_13_ARPROT;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARCACHE <= twiddle_rsc_0_13_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARBURST <= twiddle_rsc_0_13_ARBURST;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARSIZE <= twiddle_rsc_0_13_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARLEN <= twiddle_rsc_0_13_ARLEN;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_ARADDR <= twiddle_rsc_0_13_ARADDR;
  twiddle_rsc_0_13_BRESP <= peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_BRESP;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_WSTRB <= twiddle_rsc_0_13_WSTRB;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_WDATA <= twiddle_rsc_0_13_WDATA;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWREGION <= twiddle_rsc_0_13_AWREGION;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWQOS <= twiddle_rsc_0_13_AWQOS;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWPROT <= twiddle_rsc_0_13_AWPROT;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWCACHE <= twiddle_rsc_0_13_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWBURST <= twiddle_rsc_0_13_AWBURST;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWSIZE <= twiddle_rsc_0_13_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWLEN <= twiddle_rsc_0_13_AWLEN;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_AWADDR <= twiddle_rsc_0_13_AWADDR;
  peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_13_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_13_i_inst_twiddle_rsc_0_13_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_14_i_inst : peaseNTT_core_twiddle_rsc_0_14_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_14_s_tdone => twiddle_rsc_0_14_s_tdone,
      twiddle_rsc_0_14_tr_write_done => twiddle_rsc_0_14_tr_write_done,
      twiddle_rsc_0_14_RREADY => twiddle_rsc_0_14_RREADY,
      twiddle_rsc_0_14_RVALID => twiddle_rsc_0_14_RVALID,
      twiddle_rsc_0_14_RUSER => twiddle_rsc_0_14_RUSER,
      twiddle_rsc_0_14_RLAST => twiddle_rsc_0_14_RLAST,
      twiddle_rsc_0_14_RRESP => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_RRESP,
      twiddle_rsc_0_14_RDATA => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_RDATA,
      twiddle_rsc_0_14_RID => twiddle_rsc_0_14_RID,
      twiddle_rsc_0_14_ARREADY => twiddle_rsc_0_14_ARREADY,
      twiddle_rsc_0_14_ARVALID => twiddle_rsc_0_14_ARVALID,
      twiddle_rsc_0_14_ARUSER => twiddle_rsc_0_14_ARUSER,
      twiddle_rsc_0_14_ARREGION => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARREGION,
      twiddle_rsc_0_14_ARQOS => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARQOS,
      twiddle_rsc_0_14_ARPROT => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARPROT,
      twiddle_rsc_0_14_ARCACHE => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARCACHE,
      twiddle_rsc_0_14_ARLOCK => twiddle_rsc_0_14_ARLOCK,
      twiddle_rsc_0_14_ARBURST => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARBURST,
      twiddle_rsc_0_14_ARSIZE => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARSIZE,
      twiddle_rsc_0_14_ARLEN => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARLEN,
      twiddle_rsc_0_14_ARADDR => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARADDR,
      twiddle_rsc_0_14_ARID => twiddle_rsc_0_14_ARID,
      twiddle_rsc_0_14_BREADY => twiddle_rsc_0_14_BREADY,
      twiddle_rsc_0_14_BVALID => twiddle_rsc_0_14_BVALID,
      twiddle_rsc_0_14_BUSER => twiddle_rsc_0_14_BUSER,
      twiddle_rsc_0_14_BRESP => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_BRESP,
      twiddle_rsc_0_14_BID => twiddle_rsc_0_14_BID,
      twiddle_rsc_0_14_WREADY => twiddle_rsc_0_14_WREADY,
      twiddle_rsc_0_14_WVALID => twiddle_rsc_0_14_WVALID,
      twiddle_rsc_0_14_WUSER => twiddle_rsc_0_14_WUSER,
      twiddle_rsc_0_14_WLAST => twiddle_rsc_0_14_WLAST,
      twiddle_rsc_0_14_WSTRB => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_WSTRB,
      twiddle_rsc_0_14_WDATA => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_WDATA,
      twiddle_rsc_0_14_AWREADY => twiddle_rsc_0_14_AWREADY,
      twiddle_rsc_0_14_AWVALID => twiddle_rsc_0_14_AWVALID,
      twiddle_rsc_0_14_AWUSER => twiddle_rsc_0_14_AWUSER,
      twiddle_rsc_0_14_AWREGION => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWREGION,
      twiddle_rsc_0_14_AWQOS => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWQOS,
      twiddle_rsc_0_14_AWPROT => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWPROT,
      twiddle_rsc_0_14_AWCACHE => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWCACHE,
      twiddle_rsc_0_14_AWLOCK => twiddle_rsc_0_14_AWLOCK,
      twiddle_rsc_0_14_AWBURST => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWBURST,
      twiddle_rsc_0_14_AWSIZE => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWSIZE,
      twiddle_rsc_0_14_AWLEN => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWLEN,
      twiddle_rsc_0_14_AWADDR => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWADDR,
      twiddle_rsc_0_14_AWID => twiddle_rsc_0_14_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_14_i_oswt => reg_twiddle_rsc_0_6_i_oswt_cse,
      twiddle_rsc_0_14_i_wen_comp => twiddle_rsc_0_14_i_wen_comp,
      twiddle_rsc_0_14_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_i_s_raddr_core,
      twiddle_rsc_0_14_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_i_s_din_mxwt
    );
  twiddle_rsc_0_14_RRESP <= peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_RRESP;
  twiddle_rsc_0_14_RDATA <= peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_RDATA;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARREGION <= twiddle_rsc_0_14_ARREGION;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARQOS <= twiddle_rsc_0_14_ARQOS;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARPROT <= twiddle_rsc_0_14_ARPROT;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARCACHE <= twiddle_rsc_0_14_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARBURST <= twiddle_rsc_0_14_ARBURST;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARSIZE <= twiddle_rsc_0_14_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARLEN <= twiddle_rsc_0_14_ARLEN;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_ARADDR <= twiddle_rsc_0_14_ARADDR;
  twiddle_rsc_0_14_BRESP <= peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_BRESP;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_WSTRB <= twiddle_rsc_0_14_WSTRB;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_WDATA <= twiddle_rsc_0_14_WDATA;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWREGION <= twiddle_rsc_0_14_AWREGION;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWQOS <= twiddle_rsc_0_14_AWQOS;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWPROT <= twiddle_rsc_0_14_AWPROT;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWCACHE <= twiddle_rsc_0_14_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWBURST <= twiddle_rsc_0_14_AWBURST;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWSIZE <= twiddle_rsc_0_14_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWLEN <= twiddle_rsc_0_14_AWLEN;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_AWADDR <= twiddle_rsc_0_14_AWADDR;
  peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_14_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_14_i_inst_twiddle_rsc_0_14_i_s_din_mxwt;

  peaseNTT_core_twiddle_rsc_0_15_i_inst : peaseNTT_core_twiddle_rsc_0_15_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_rsc_0_15_s_tdone => twiddle_rsc_0_15_s_tdone,
      twiddle_rsc_0_15_tr_write_done => twiddle_rsc_0_15_tr_write_done,
      twiddle_rsc_0_15_RREADY => twiddle_rsc_0_15_RREADY,
      twiddle_rsc_0_15_RVALID => twiddle_rsc_0_15_RVALID,
      twiddle_rsc_0_15_RUSER => twiddle_rsc_0_15_RUSER,
      twiddle_rsc_0_15_RLAST => twiddle_rsc_0_15_RLAST,
      twiddle_rsc_0_15_RRESP => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_RRESP,
      twiddle_rsc_0_15_RDATA => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_RDATA,
      twiddle_rsc_0_15_RID => twiddle_rsc_0_15_RID,
      twiddle_rsc_0_15_ARREADY => twiddle_rsc_0_15_ARREADY,
      twiddle_rsc_0_15_ARVALID => twiddle_rsc_0_15_ARVALID,
      twiddle_rsc_0_15_ARUSER => twiddle_rsc_0_15_ARUSER,
      twiddle_rsc_0_15_ARREGION => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARREGION,
      twiddle_rsc_0_15_ARQOS => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARQOS,
      twiddle_rsc_0_15_ARPROT => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARPROT,
      twiddle_rsc_0_15_ARCACHE => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARCACHE,
      twiddle_rsc_0_15_ARLOCK => twiddle_rsc_0_15_ARLOCK,
      twiddle_rsc_0_15_ARBURST => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARBURST,
      twiddle_rsc_0_15_ARSIZE => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARSIZE,
      twiddle_rsc_0_15_ARLEN => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARLEN,
      twiddle_rsc_0_15_ARADDR => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARADDR,
      twiddle_rsc_0_15_ARID => twiddle_rsc_0_15_ARID,
      twiddle_rsc_0_15_BREADY => twiddle_rsc_0_15_BREADY,
      twiddle_rsc_0_15_BVALID => twiddle_rsc_0_15_BVALID,
      twiddle_rsc_0_15_BUSER => twiddle_rsc_0_15_BUSER,
      twiddle_rsc_0_15_BRESP => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_BRESP,
      twiddle_rsc_0_15_BID => twiddle_rsc_0_15_BID,
      twiddle_rsc_0_15_WREADY => twiddle_rsc_0_15_WREADY,
      twiddle_rsc_0_15_WVALID => twiddle_rsc_0_15_WVALID,
      twiddle_rsc_0_15_WUSER => twiddle_rsc_0_15_WUSER,
      twiddle_rsc_0_15_WLAST => twiddle_rsc_0_15_WLAST,
      twiddle_rsc_0_15_WSTRB => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_WSTRB,
      twiddle_rsc_0_15_WDATA => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_WDATA,
      twiddle_rsc_0_15_AWREADY => twiddle_rsc_0_15_AWREADY,
      twiddle_rsc_0_15_AWVALID => twiddle_rsc_0_15_AWVALID,
      twiddle_rsc_0_15_AWUSER => twiddle_rsc_0_15_AWUSER,
      twiddle_rsc_0_15_AWREGION => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWREGION,
      twiddle_rsc_0_15_AWQOS => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWQOS,
      twiddle_rsc_0_15_AWPROT => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWPROT,
      twiddle_rsc_0_15_AWCACHE => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWCACHE,
      twiddle_rsc_0_15_AWLOCK => twiddle_rsc_0_15_AWLOCK,
      twiddle_rsc_0_15_AWBURST => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWBURST,
      twiddle_rsc_0_15_AWSIZE => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWSIZE,
      twiddle_rsc_0_15_AWLEN => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWLEN,
      twiddle_rsc_0_15_AWADDR => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWADDR,
      twiddle_rsc_0_15_AWID => twiddle_rsc_0_15_AWID,
      core_wen => core_wen,
      twiddle_rsc_0_15_i_oswt => reg_twiddle_rsc_0_7_i_oswt_cse,
      twiddle_rsc_0_15_i_wen_comp => twiddle_rsc_0_15_i_wen_comp,
      twiddle_rsc_0_15_i_s_raddr_core => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_i_s_raddr_core,
      twiddle_rsc_0_15_i_s_din_mxwt => peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_i_s_din_mxwt
    );
  twiddle_rsc_0_15_RRESP <= peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_RRESP;
  twiddle_rsc_0_15_RDATA <= peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_RDATA;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARREGION <= twiddle_rsc_0_15_ARREGION;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARQOS <= twiddle_rsc_0_15_ARQOS;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARPROT <= twiddle_rsc_0_15_ARPROT;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARCACHE <= twiddle_rsc_0_15_ARCACHE;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARBURST <= twiddle_rsc_0_15_ARBURST;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARSIZE <= twiddle_rsc_0_15_ARSIZE;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARLEN <= twiddle_rsc_0_15_ARLEN;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_ARADDR <= twiddle_rsc_0_15_ARADDR;
  twiddle_rsc_0_15_BRESP <= peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_BRESP;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_WSTRB <= twiddle_rsc_0_15_WSTRB;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_WDATA <= twiddle_rsc_0_15_WDATA;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWREGION <= twiddle_rsc_0_15_AWREGION;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWQOS <= twiddle_rsc_0_15_AWQOS;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWPROT <= twiddle_rsc_0_15_AWPROT;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWCACHE <= twiddle_rsc_0_15_AWCACHE;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWBURST <= twiddle_rsc_0_15_AWBURST;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWSIZE <= twiddle_rsc_0_15_AWSIZE;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWLEN <= twiddle_rsc_0_15_AWLEN;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_AWADDR <= twiddle_rsc_0_15_AWADDR;
  peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_rsc_0_15_i_s_din_mxwt <= peaseNTT_core_twiddle_rsc_0_15_i_inst_twiddle_rsc_0_15_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_0_i_inst : peaseNTT_core_twiddle_h_rsc_0_0_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_0_s_tdone => twiddle_h_rsc_0_0_s_tdone,
      twiddle_h_rsc_0_0_tr_write_done => twiddle_h_rsc_0_0_tr_write_done,
      twiddle_h_rsc_0_0_RREADY => twiddle_h_rsc_0_0_RREADY,
      twiddle_h_rsc_0_0_RVALID => twiddle_h_rsc_0_0_RVALID,
      twiddle_h_rsc_0_0_RUSER => twiddle_h_rsc_0_0_RUSER,
      twiddle_h_rsc_0_0_RLAST => twiddle_h_rsc_0_0_RLAST,
      twiddle_h_rsc_0_0_RRESP => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_RRESP,
      twiddle_h_rsc_0_0_RDATA => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_RDATA,
      twiddle_h_rsc_0_0_RID => twiddle_h_rsc_0_0_RID,
      twiddle_h_rsc_0_0_ARREADY => twiddle_h_rsc_0_0_ARREADY,
      twiddle_h_rsc_0_0_ARVALID => twiddle_h_rsc_0_0_ARVALID,
      twiddle_h_rsc_0_0_ARUSER => twiddle_h_rsc_0_0_ARUSER,
      twiddle_h_rsc_0_0_ARREGION => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARREGION,
      twiddle_h_rsc_0_0_ARQOS => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARQOS,
      twiddle_h_rsc_0_0_ARPROT => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARPROT,
      twiddle_h_rsc_0_0_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARCACHE,
      twiddle_h_rsc_0_0_ARLOCK => twiddle_h_rsc_0_0_ARLOCK,
      twiddle_h_rsc_0_0_ARBURST => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARBURST,
      twiddle_h_rsc_0_0_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARSIZE,
      twiddle_h_rsc_0_0_ARLEN => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARLEN,
      twiddle_h_rsc_0_0_ARADDR => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARADDR,
      twiddle_h_rsc_0_0_ARID => twiddle_h_rsc_0_0_ARID,
      twiddle_h_rsc_0_0_BREADY => twiddle_h_rsc_0_0_BREADY,
      twiddle_h_rsc_0_0_BVALID => twiddle_h_rsc_0_0_BVALID,
      twiddle_h_rsc_0_0_BUSER => twiddle_h_rsc_0_0_BUSER,
      twiddle_h_rsc_0_0_BRESP => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_BRESP,
      twiddle_h_rsc_0_0_BID => twiddle_h_rsc_0_0_BID,
      twiddle_h_rsc_0_0_WREADY => twiddle_h_rsc_0_0_WREADY,
      twiddle_h_rsc_0_0_WVALID => twiddle_h_rsc_0_0_WVALID,
      twiddle_h_rsc_0_0_WUSER => twiddle_h_rsc_0_0_WUSER,
      twiddle_h_rsc_0_0_WLAST => twiddle_h_rsc_0_0_WLAST,
      twiddle_h_rsc_0_0_WSTRB => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_WSTRB,
      twiddle_h_rsc_0_0_WDATA => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_WDATA,
      twiddle_h_rsc_0_0_AWREADY => twiddle_h_rsc_0_0_AWREADY,
      twiddle_h_rsc_0_0_AWVALID => twiddle_h_rsc_0_0_AWVALID,
      twiddle_h_rsc_0_0_AWUSER => twiddle_h_rsc_0_0_AWUSER,
      twiddle_h_rsc_0_0_AWREGION => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWREGION,
      twiddle_h_rsc_0_0_AWQOS => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWQOS,
      twiddle_h_rsc_0_0_AWPROT => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWPROT,
      twiddle_h_rsc_0_0_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWCACHE,
      twiddle_h_rsc_0_0_AWLOCK => twiddle_h_rsc_0_0_AWLOCK,
      twiddle_h_rsc_0_0_AWBURST => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWBURST,
      twiddle_h_rsc_0_0_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWSIZE,
      twiddle_h_rsc_0_0_AWLEN => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWLEN,
      twiddle_h_rsc_0_0_AWADDR => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWADDR,
      twiddle_h_rsc_0_0_AWID => twiddle_h_rsc_0_0_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_0_i_oswt => reg_twiddle_rsc_0_0_i_oswt_cse,
      twiddle_h_rsc_0_0_i_wen_comp => twiddle_h_rsc_0_0_i_wen_comp,
      twiddle_h_rsc_0_0_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_i_s_raddr_core,
      twiddle_h_rsc_0_0_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_i_s_din_mxwt
    );
  twiddle_h_rsc_0_0_RRESP <= peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_RRESP;
  twiddle_h_rsc_0_0_RDATA <= peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARREGION <= twiddle_h_rsc_0_0_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARQOS <= twiddle_h_rsc_0_0_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARPROT <= twiddle_h_rsc_0_0_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARCACHE <= twiddle_h_rsc_0_0_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARBURST <= twiddle_h_rsc_0_0_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARSIZE <= twiddle_h_rsc_0_0_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARLEN <= twiddle_h_rsc_0_0_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_ARADDR <= twiddle_h_rsc_0_0_ARADDR;
  twiddle_h_rsc_0_0_BRESP <= peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_WSTRB <= twiddle_h_rsc_0_0_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_WDATA <= twiddle_h_rsc_0_0_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWREGION <= twiddle_h_rsc_0_0_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWQOS <= twiddle_h_rsc_0_0_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWPROT <= twiddle_h_rsc_0_0_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWCACHE <= twiddle_h_rsc_0_0_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWBURST <= twiddle_h_rsc_0_0_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWSIZE <= twiddle_h_rsc_0_0_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWLEN <= twiddle_h_rsc_0_0_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_AWADDR <= twiddle_h_rsc_0_0_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_i_s_raddr_core <= '0'
      & twiddle_h_rsc_0_0_i_s_raddr_core_4 & reg_twiddle_rsc_0_0_i_s_raddr_core_3_0_cse;
  twiddle_h_rsc_0_0_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_0_i_inst_twiddle_h_rsc_0_0_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_1_i_inst : peaseNTT_core_twiddle_h_rsc_0_1_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_1_s_tdone => twiddle_h_rsc_0_1_s_tdone,
      twiddle_h_rsc_0_1_tr_write_done => twiddle_h_rsc_0_1_tr_write_done,
      twiddle_h_rsc_0_1_RREADY => twiddle_h_rsc_0_1_RREADY,
      twiddle_h_rsc_0_1_RVALID => twiddle_h_rsc_0_1_RVALID,
      twiddle_h_rsc_0_1_RUSER => twiddle_h_rsc_0_1_RUSER,
      twiddle_h_rsc_0_1_RLAST => twiddle_h_rsc_0_1_RLAST,
      twiddle_h_rsc_0_1_RRESP => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_RRESP,
      twiddle_h_rsc_0_1_RDATA => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_RDATA,
      twiddle_h_rsc_0_1_RID => twiddle_h_rsc_0_1_RID,
      twiddle_h_rsc_0_1_ARREADY => twiddle_h_rsc_0_1_ARREADY,
      twiddle_h_rsc_0_1_ARVALID => twiddle_h_rsc_0_1_ARVALID,
      twiddle_h_rsc_0_1_ARUSER => twiddle_h_rsc_0_1_ARUSER,
      twiddle_h_rsc_0_1_ARREGION => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARREGION,
      twiddle_h_rsc_0_1_ARQOS => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARQOS,
      twiddle_h_rsc_0_1_ARPROT => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARPROT,
      twiddle_h_rsc_0_1_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARCACHE,
      twiddle_h_rsc_0_1_ARLOCK => twiddle_h_rsc_0_1_ARLOCK,
      twiddle_h_rsc_0_1_ARBURST => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARBURST,
      twiddle_h_rsc_0_1_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARSIZE,
      twiddle_h_rsc_0_1_ARLEN => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARLEN,
      twiddle_h_rsc_0_1_ARADDR => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARADDR,
      twiddle_h_rsc_0_1_ARID => twiddle_h_rsc_0_1_ARID,
      twiddle_h_rsc_0_1_BREADY => twiddle_h_rsc_0_1_BREADY,
      twiddle_h_rsc_0_1_BVALID => twiddle_h_rsc_0_1_BVALID,
      twiddle_h_rsc_0_1_BUSER => twiddle_h_rsc_0_1_BUSER,
      twiddle_h_rsc_0_1_BRESP => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_BRESP,
      twiddle_h_rsc_0_1_BID => twiddle_h_rsc_0_1_BID,
      twiddle_h_rsc_0_1_WREADY => twiddle_h_rsc_0_1_WREADY,
      twiddle_h_rsc_0_1_WVALID => twiddle_h_rsc_0_1_WVALID,
      twiddle_h_rsc_0_1_WUSER => twiddle_h_rsc_0_1_WUSER,
      twiddle_h_rsc_0_1_WLAST => twiddle_h_rsc_0_1_WLAST,
      twiddle_h_rsc_0_1_WSTRB => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_WSTRB,
      twiddle_h_rsc_0_1_WDATA => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_WDATA,
      twiddle_h_rsc_0_1_AWREADY => twiddle_h_rsc_0_1_AWREADY,
      twiddle_h_rsc_0_1_AWVALID => twiddle_h_rsc_0_1_AWVALID,
      twiddle_h_rsc_0_1_AWUSER => twiddle_h_rsc_0_1_AWUSER,
      twiddle_h_rsc_0_1_AWREGION => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWREGION,
      twiddle_h_rsc_0_1_AWQOS => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWQOS,
      twiddle_h_rsc_0_1_AWPROT => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWPROT,
      twiddle_h_rsc_0_1_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWCACHE,
      twiddle_h_rsc_0_1_AWLOCK => twiddle_h_rsc_0_1_AWLOCK,
      twiddle_h_rsc_0_1_AWBURST => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWBURST,
      twiddle_h_rsc_0_1_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWSIZE,
      twiddle_h_rsc_0_1_AWLEN => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWLEN,
      twiddle_h_rsc_0_1_AWADDR => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWADDR,
      twiddle_h_rsc_0_1_AWID => twiddle_h_rsc_0_1_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_1_i_oswt => reg_twiddle_rsc_0_1_i_oswt_cse,
      twiddle_h_rsc_0_1_i_wen_comp => twiddle_h_rsc_0_1_i_wen_comp,
      twiddle_h_rsc_0_1_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_i_s_raddr_core,
      twiddle_h_rsc_0_1_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_i_s_din_mxwt
    );
  twiddle_h_rsc_0_1_RRESP <= peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_RRESP;
  twiddle_h_rsc_0_1_RDATA <= peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARREGION <= twiddle_h_rsc_0_1_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARQOS <= twiddle_h_rsc_0_1_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARPROT <= twiddle_h_rsc_0_1_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARCACHE <= twiddle_h_rsc_0_1_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARBURST <= twiddle_h_rsc_0_1_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARSIZE <= twiddle_h_rsc_0_1_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARLEN <= twiddle_h_rsc_0_1_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_ARADDR <= twiddle_h_rsc_0_1_ARADDR;
  twiddle_h_rsc_0_1_BRESP <= peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_WSTRB <= twiddle_h_rsc_0_1_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_WDATA <= twiddle_h_rsc_0_1_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWREGION <= twiddle_h_rsc_0_1_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWQOS <= twiddle_h_rsc_0_1_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWPROT <= twiddle_h_rsc_0_1_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWCACHE <= twiddle_h_rsc_0_1_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWBURST <= twiddle_h_rsc_0_1_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWSIZE <= twiddle_h_rsc_0_1_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWLEN <= twiddle_h_rsc_0_1_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_AWADDR <= twiddle_h_rsc_0_1_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_1_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_1_i_inst_twiddle_h_rsc_0_1_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_2_i_inst : peaseNTT_core_twiddle_h_rsc_0_2_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_2_s_tdone => twiddle_h_rsc_0_2_s_tdone,
      twiddle_h_rsc_0_2_tr_write_done => twiddle_h_rsc_0_2_tr_write_done,
      twiddle_h_rsc_0_2_RREADY => twiddle_h_rsc_0_2_RREADY,
      twiddle_h_rsc_0_2_RVALID => twiddle_h_rsc_0_2_RVALID,
      twiddle_h_rsc_0_2_RUSER => twiddle_h_rsc_0_2_RUSER,
      twiddle_h_rsc_0_2_RLAST => twiddle_h_rsc_0_2_RLAST,
      twiddle_h_rsc_0_2_RRESP => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_RRESP,
      twiddle_h_rsc_0_2_RDATA => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_RDATA,
      twiddle_h_rsc_0_2_RID => twiddle_h_rsc_0_2_RID,
      twiddle_h_rsc_0_2_ARREADY => twiddle_h_rsc_0_2_ARREADY,
      twiddle_h_rsc_0_2_ARVALID => twiddle_h_rsc_0_2_ARVALID,
      twiddle_h_rsc_0_2_ARUSER => twiddle_h_rsc_0_2_ARUSER,
      twiddle_h_rsc_0_2_ARREGION => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARREGION,
      twiddle_h_rsc_0_2_ARQOS => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARQOS,
      twiddle_h_rsc_0_2_ARPROT => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARPROT,
      twiddle_h_rsc_0_2_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARCACHE,
      twiddle_h_rsc_0_2_ARLOCK => twiddle_h_rsc_0_2_ARLOCK,
      twiddle_h_rsc_0_2_ARBURST => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARBURST,
      twiddle_h_rsc_0_2_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARSIZE,
      twiddle_h_rsc_0_2_ARLEN => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARLEN,
      twiddle_h_rsc_0_2_ARADDR => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARADDR,
      twiddle_h_rsc_0_2_ARID => twiddle_h_rsc_0_2_ARID,
      twiddle_h_rsc_0_2_BREADY => twiddle_h_rsc_0_2_BREADY,
      twiddle_h_rsc_0_2_BVALID => twiddle_h_rsc_0_2_BVALID,
      twiddle_h_rsc_0_2_BUSER => twiddle_h_rsc_0_2_BUSER,
      twiddle_h_rsc_0_2_BRESP => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_BRESP,
      twiddle_h_rsc_0_2_BID => twiddle_h_rsc_0_2_BID,
      twiddle_h_rsc_0_2_WREADY => twiddle_h_rsc_0_2_WREADY,
      twiddle_h_rsc_0_2_WVALID => twiddle_h_rsc_0_2_WVALID,
      twiddle_h_rsc_0_2_WUSER => twiddle_h_rsc_0_2_WUSER,
      twiddle_h_rsc_0_2_WLAST => twiddle_h_rsc_0_2_WLAST,
      twiddle_h_rsc_0_2_WSTRB => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_WSTRB,
      twiddle_h_rsc_0_2_WDATA => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_WDATA,
      twiddle_h_rsc_0_2_AWREADY => twiddle_h_rsc_0_2_AWREADY,
      twiddle_h_rsc_0_2_AWVALID => twiddle_h_rsc_0_2_AWVALID,
      twiddle_h_rsc_0_2_AWUSER => twiddle_h_rsc_0_2_AWUSER,
      twiddle_h_rsc_0_2_AWREGION => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWREGION,
      twiddle_h_rsc_0_2_AWQOS => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWQOS,
      twiddle_h_rsc_0_2_AWPROT => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWPROT,
      twiddle_h_rsc_0_2_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWCACHE,
      twiddle_h_rsc_0_2_AWLOCK => twiddle_h_rsc_0_2_AWLOCK,
      twiddle_h_rsc_0_2_AWBURST => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWBURST,
      twiddle_h_rsc_0_2_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWSIZE,
      twiddle_h_rsc_0_2_AWLEN => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWLEN,
      twiddle_h_rsc_0_2_AWADDR => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWADDR,
      twiddle_h_rsc_0_2_AWID => twiddle_h_rsc_0_2_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_2_i_oswt => reg_twiddle_rsc_0_2_i_oswt_cse,
      twiddle_h_rsc_0_2_i_wen_comp => twiddle_h_rsc_0_2_i_wen_comp,
      twiddle_h_rsc_0_2_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_i_s_raddr_core,
      twiddle_h_rsc_0_2_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_i_s_din_mxwt
    );
  twiddle_h_rsc_0_2_RRESP <= peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_RRESP;
  twiddle_h_rsc_0_2_RDATA <= peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARREGION <= twiddle_h_rsc_0_2_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARQOS <= twiddle_h_rsc_0_2_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARPROT <= twiddle_h_rsc_0_2_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARCACHE <= twiddle_h_rsc_0_2_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARBURST <= twiddle_h_rsc_0_2_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARSIZE <= twiddle_h_rsc_0_2_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARLEN <= twiddle_h_rsc_0_2_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_ARADDR <= twiddle_h_rsc_0_2_ARADDR;
  twiddle_h_rsc_0_2_BRESP <= peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_WSTRB <= twiddle_h_rsc_0_2_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_WDATA <= twiddle_h_rsc_0_2_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWREGION <= twiddle_h_rsc_0_2_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWQOS <= twiddle_h_rsc_0_2_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWPROT <= twiddle_h_rsc_0_2_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWCACHE <= twiddle_h_rsc_0_2_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWBURST <= twiddle_h_rsc_0_2_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWSIZE <= twiddle_h_rsc_0_2_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWLEN <= twiddle_h_rsc_0_2_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_AWADDR <= twiddle_h_rsc_0_2_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_2_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_2_i_inst_twiddle_h_rsc_0_2_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_3_i_inst : peaseNTT_core_twiddle_h_rsc_0_3_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_3_s_tdone => twiddle_h_rsc_0_3_s_tdone,
      twiddle_h_rsc_0_3_tr_write_done => twiddle_h_rsc_0_3_tr_write_done,
      twiddle_h_rsc_0_3_RREADY => twiddle_h_rsc_0_3_RREADY,
      twiddle_h_rsc_0_3_RVALID => twiddle_h_rsc_0_3_RVALID,
      twiddle_h_rsc_0_3_RUSER => twiddle_h_rsc_0_3_RUSER,
      twiddle_h_rsc_0_3_RLAST => twiddle_h_rsc_0_3_RLAST,
      twiddle_h_rsc_0_3_RRESP => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_RRESP,
      twiddle_h_rsc_0_3_RDATA => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_RDATA,
      twiddle_h_rsc_0_3_RID => twiddle_h_rsc_0_3_RID,
      twiddle_h_rsc_0_3_ARREADY => twiddle_h_rsc_0_3_ARREADY,
      twiddle_h_rsc_0_3_ARVALID => twiddle_h_rsc_0_3_ARVALID,
      twiddle_h_rsc_0_3_ARUSER => twiddle_h_rsc_0_3_ARUSER,
      twiddle_h_rsc_0_3_ARREGION => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARREGION,
      twiddle_h_rsc_0_3_ARQOS => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARQOS,
      twiddle_h_rsc_0_3_ARPROT => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARPROT,
      twiddle_h_rsc_0_3_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARCACHE,
      twiddle_h_rsc_0_3_ARLOCK => twiddle_h_rsc_0_3_ARLOCK,
      twiddle_h_rsc_0_3_ARBURST => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARBURST,
      twiddle_h_rsc_0_3_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARSIZE,
      twiddle_h_rsc_0_3_ARLEN => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARLEN,
      twiddle_h_rsc_0_3_ARADDR => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARADDR,
      twiddle_h_rsc_0_3_ARID => twiddle_h_rsc_0_3_ARID,
      twiddle_h_rsc_0_3_BREADY => twiddle_h_rsc_0_3_BREADY,
      twiddle_h_rsc_0_3_BVALID => twiddle_h_rsc_0_3_BVALID,
      twiddle_h_rsc_0_3_BUSER => twiddle_h_rsc_0_3_BUSER,
      twiddle_h_rsc_0_3_BRESP => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_BRESP,
      twiddle_h_rsc_0_3_BID => twiddle_h_rsc_0_3_BID,
      twiddle_h_rsc_0_3_WREADY => twiddle_h_rsc_0_3_WREADY,
      twiddle_h_rsc_0_3_WVALID => twiddle_h_rsc_0_3_WVALID,
      twiddle_h_rsc_0_3_WUSER => twiddle_h_rsc_0_3_WUSER,
      twiddle_h_rsc_0_3_WLAST => twiddle_h_rsc_0_3_WLAST,
      twiddle_h_rsc_0_3_WSTRB => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_WSTRB,
      twiddle_h_rsc_0_3_WDATA => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_WDATA,
      twiddle_h_rsc_0_3_AWREADY => twiddle_h_rsc_0_3_AWREADY,
      twiddle_h_rsc_0_3_AWVALID => twiddle_h_rsc_0_3_AWVALID,
      twiddle_h_rsc_0_3_AWUSER => twiddle_h_rsc_0_3_AWUSER,
      twiddle_h_rsc_0_3_AWREGION => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWREGION,
      twiddle_h_rsc_0_3_AWQOS => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWQOS,
      twiddle_h_rsc_0_3_AWPROT => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWPROT,
      twiddle_h_rsc_0_3_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWCACHE,
      twiddle_h_rsc_0_3_AWLOCK => twiddle_h_rsc_0_3_AWLOCK,
      twiddle_h_rsc_0_3_AWBURST => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWBURST,
      twiddle_h_rsc_0_3_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWSIZE,
      twiddle_h_rsc_0_3_AWLEN => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWLEN,
      twiddle_h_rsc_0_3_AWADDR => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWADDR,
      twiddle_h_rsc_0_3_AWID => twiddle_h_rsc_0_3_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_3_i_oswt => reg_twiddle_rsc_0_3_i_oswt_cse,
      twiddle_h_rsc_0_3_i_wen_comp => twiddle_h_rsc_0_3_i_wen_comp,
      twiddle_h_rsc_0_3_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_i_s_raddr_core,
      twiddle_h_rsc_0_3_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_i_s_din_mxwt
    );
  twiddle_h_rsc_0_3_RRESP <= peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_RRESP;
  twiddle_h_rsc_0_3_RDATA <= peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARREGION <= twiddle_h_rsc_0_3_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARQOS <= twiddle_h_rsc_0_3_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARPROT <= twiddle_h_rsc_0_3_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARCACHE <= twiddle_h_rsc_0_3_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARBURST <= twiddle_h_rsc_0_3_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARSIZE <= twiddle_h_rsc_0_3_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARLEN <= twiddle_h_rsc_0_3_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_ARADDR <= twiddle_h_rsc_0_3_ARADDR;
  twiddle_h_rsc_0_3_BRESP <= peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_WSTRB <= twiddle_h_rsc_0_3_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_WDATA <= twiddle_h_rsc_0_3_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWREGION <= twiddle_h_rsc_0_3_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWQOS <= twiddle_h_rsc_0_3_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWPROT <= twiddle_h_rsc_0_3_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWCACHE <= twiddle_h_rsc_0_3_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWBURST <= twiddle_h_rsc_0_3_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWSIZE <= twiddle_h_rsc_0_3_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWLEN <= twiddle_h_rsc_0_3_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_AWADDR <= twiddle_h_rsc_0_3_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_3_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_3_i_inst_twiddle_h_rsc_0_3_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_4_i_inst : peaseNTT_core_twiddle_h_rsc_0_4_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_4_s_tdone => twiddle_h_rsc_0_4_s_tdone,
      twiddle_h_rsc_0_4_tr_write_done => twiddle_h_rsc_0_4_tr_write_done,
      twiddle_h_rsc_0_4_RREADY => twiddle_h_rsc_0_4_RREADY,
      twiddle_h_rsc_0_4_RVALID => twiddle_h_rsc_0_4_RVALID,
      twiddle_h_rsc_0_4_RUSER => twiddle_h_rsc_0_4_RUSER,
      twiddle_h_rsc_0_4_RLAST => twiddle_h_rsc_0_4_RLAST,
      twiddle_h_rsc_0_4_RRESP => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_RRESP,
      twiddle_h_rsc_0_4_RDATA => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_RDATA,
      twiddle_h_rsc_0_4_RID => twiddle_h_rsc_0_4_RID,
      twiddle_h_rsc_0_4_ARREADY => twiddle_h_rsc_0_4_ARREADY,
      twiddle_h_rsc_0_4_ARVALID => twiddle_h_rsc_0_4_ARVALID,
      twiddle_h_rsc_0_4_ARUSER => twiddle_h_rsc_0_4_ARUSER,
      twiddle_h_rsc_0_4_ARREGION => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARREGION,
      twiddle_h_rsc_0_4_ARQOS => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARQOS,
      twiddle_h_rsc_0_4_ARPROT => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARPROT,
      twiddle_h_rsc_0_4_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARCACHE,
      twiddle_h_rsc_0_4_ARLOCK => twiddle_h_rsc_0_4_ARLOCK,
      twiddle_h_rsc_0_4_ARBURST => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARBURST,
      twiddle_h_rsc_0_4_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARSIZE,
      twiddle_h_rsc_0_4_ARLEN => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARLEN,
      twiddle_h_rsc_0_4_ARADDR => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARADDR,
      twiddle_h_rsc_0_4_ARID => twiddle_h_rsc_0_4_ARID,
      twiddle_h_rsc_0_4_BREADY => twiddle_h_rsc_0_4_BREADY,
      twiddle_h_rsc_0_4_BVALID => twiddle_h_rsc_0_4_BVALID,
      twiddle_h_rsc_0_4_BUSER => twiddle_h_rsc_0_4_BUSER,
      twiddle_h_rsc_0_4_BRESP => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_BRESP,
      twiddle_h_rsc_0_4_BID => twiddle_h_rsc_0_4_BID,
      twiddle_h_rsc_0_4_WREADY => twiddle_h_rsc_0_4_WREADY,
      twiddle_h_rsc_0_4_WVALID => twiddle_h_rsc_0_4_WVALID,
      twiddle_h_rsc_0_4_WUSER => twiddle_h_rsc_0_4_WUSER,
      twiddle_h_rsc_0_4_WLAST => twiddle_h_rsc_0_4_WLAST,
      twiddle_h_rsc_0_4_WSTRB => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_WSTRB,
      twiddle_h_rsc_0_4_WDATA => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_WDATA,
      twiddle_h_rsc_0_4_AWREADY => twiddle_h_rsc_0_4_AWREADY,
      twiddle_h_rsc_0_4_AWVALID => twiddle_h_rsc_0_4_AWVALID,
      twiddle_h_rsc_0_4_AWUSER => twiddle_h_rsc_0_4_AWUSER,
      twiddle_h_rsc_0_4_AWREGION => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWREGION,
      twiddle_h_rsc_0_4_AWQOS => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWQOS,
      twiddle_h_rsc_0_4_AWPROT => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWPROT,
      twiddle_h_rsc_0_4_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWCACHE,
      twiddle_h_rsc_0_4_AWLOCK => twiddle_h_rsc_0_4_AWLOCK,
      twiddle_h_rsc_0_4_AWBURST => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWBURST,
      twiddle_h_rsc_0_4_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWSIZE,
      twiddle_h_rsc_0_4_AWLEN => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWLEN,
      twiddle_h_rsc_0_4_AWADDR => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWADDR,
      twiddle_h_rsc_0_4_AWID => twiddle_h_rsc_0_4_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_4_i_oswt => reg_twiddle_rsc_0_4_i_oswt_cse,
      twiddle_h_rsc_0_4_i_wen_comp => twiddle_h_rsc_0_4_i_wen_comp,
      twiddle_h_rsc_0_4_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_i_s_raddr_core,
      twiddle_h_rsc_0_4_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_i_s_din_mxwt
    );
  twiddle_h_rsc_0_4_RRESP <= peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_RRESP;
  twiddle_h_rsc_0_4_RDATA <= peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARREGION <= twiddle_h_rsc_0_4_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARQOS <= twiddle_h_rsc_0_4_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARPROT <= twiddle_h_rsc_0_4_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARCACHE <= twiddle_h_rsc_0_4_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARBURST <= twiddle_h_rsc_0_4_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARSIZE <= twiddle_h_rsc_0_4_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARLEN <= twiddle_h_rsc_0_4_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_ARADDR <= twiddle_h_rsc_0_4_ARADDR;
  twiddle_h_rsc_0_4_BRESP <= peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_WSTRB <= twiddle_h_rsc_0_4_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_WDATA <= twiddle_h_rsc_0_4_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWREGION <= twiddle_h_rsc_0_4_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWQOS <= twiddle_h_rsc_0_4_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWPROT <= twiddle_h_rsc_0_4_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWCACHE <= twiddle_h_rsc_0_4_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWBURST <= twiddle_h_rsc_0_4_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWSIZE <= twiddle_h_rsc_0_4_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWLEN <= twiddle_h_rsc_0_4_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_AWADDR <= twiddle_h_rsc_0_4_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_4_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_4_i_inst_twiddle_h_rsc_0_4_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_5_i_inst : peaseNTT_core_twiddle_h_rsc_0_5_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_5_s_tdone => twiddle_h_rsc_0_5_s_tdone,
      twiddle_h_rsc_0_5_tr_write_done => twiddle_h_rsc_0_5_tr_write_done,
      twiddle_h_rsc_0_5_RREADY => twiddle_h_rsc_0_5_RREADY,
      twiddle_h_rsc_0_5_RVALID => twiddle_h_rsc_0_5_RVALID,
      twiddle_h_rsc_0_5_RUSER => twiddle_h_rsc_0_5_RUSER,
      twiddle_h_rsc_0_5_RLAST => twiddle_h_rsc_0_5_RLAST,
      twiddle_h_rsc_0_5_RRESP => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_RRESP,
      twiddle_h_rsc_0_5_RDATA => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_RDATA,
      twiddle_h_rsc_0_5_RID => twiddle_h_rsc_0_5_RID,
      twiddle_h_rsc_0_5_ARREADY => twiddle_h_rsc_0_5_ARREADY,
      twiddle_h_rsc_0_5_ARVALID => twiddle_h_rsc_0_5_ARVALID,
      twiddle_h_rsc_0_5_ARUSER => twiddle_h_rsc_0_5_ARUSER,
      twiddle_h_rsc_0_5_ARREGION => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARREGION,
      twiddle_h_rsc_0_5_ARQOS => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARQOS,
      twiddle_h_rsc_0_5_ARPROT => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARPROT,
      twiddle_h_rsc_0_5_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARCACHE,
      twiddle_h_rsc_0_5_ARLOCK => twiddle_h_rsc_0_5_ARLOCK,
      twiddle_h_rsc_0_5_ARBURST => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARBURST,
      twiddle_h_rsc_0_5_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARSIZE,
      twiddle_h_rsc_0_5_ARLEN => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARLEN,
      twiddle_h_rsc_0_5_ARADDR => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARADDR,
      twiddle_h_rsc_0_5_ARID => twiddle_h_rsc_0_5_ARID,
      twiddle_h_rsc_0_5_BREADY => twiddle_h_rsc_0_5_BREADY,
      twiddle_h_rsc_0_5_BVALID => twiddle_h_rsc_0_5_BVALID,
      twiddle_h_rsc_0_5_BUSER => twiddle_h_rsc_0_5_BUSER,
      twiddle_h_rsc_0_5_BRESP => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_BRESP,
      twiddle_h_rsc_0_5_BID => twiddle_h_rsc_0_5_BID,
      twiddle_h_rsc_0_5_WREADY => twiddle_h_rsc_0_5_WREADY,
      twiddle_h_rsc_0_5_WVALID => twiddle_h_rsc_0_5_WVALID,
      twiddle_h_rsc_0_5_WUSER => twiddle_h_rsc_0_5_WUSER,
      twiddle_h_rsc_0_5_WLAST => twiddle_h_rsc_0_5_WLAST,
      twiddle_h_rsc_0_5_WSTRB => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_WSTRB,
      twiddle_h_rsc_0_5_WDATA => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_WDATA,
      twiddle_h_rsc_0_5_AWREADY => twiddle_h_rsc_0_5_AWREADY,
      twiddle_h_rsc_0_5_AWVALID => twiddle_h_rsc_0_5_AWVALID,
      twiddle_h_rsc_0_5_AWUSER => twiddle_h_rsc_0_5_AWUSER,
      twiddle_h_rsc_0_5_AWREGION => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWREGION,
      twiddle_h_rsc_0_5_AWQOS => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWQOS,
      twiddle_h_rsc_0_5_AWPROT => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWPROT,
      twiddle_h_rsc_0_5_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWCACHE,
      twiddle_h_rsc_0_5_AWLOCK => twiddle_h_rsc_0_5_AWLOCK,
      twiddle_h_rsc_0_5_AWBURST => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWBURST,
      twiddle_h_rsc_0_5_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWSIZE,
      twiddle_h_rsc_0_5_AWLEN => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWLEN,
      twiddle_h_rsc_0_5_AWADDR => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWADDR,
      twiddle_h_rsc_0_5_AWID => twiddle_h_rsc_0_5_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_5_i_oswt => reg_twiddle_rsc_0_5_i_oswt_cse,
      twiddle_h_rsc_0_5_i_wen_comp => twiddle_h_rsc_0_5_i_wen_comp,
      twiddle_h_rsc_0_5_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_i_s_raddr_core,
      twiddle_h_rsc_0_5_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_i_s_din_mxwt
    );
  twiddle_h_rsc_0_5_RRESP <= peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_RRESP;
  twiddle_h_rsc_0_5_RDATA <= peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARREGION <= twiddle_h_rsc_0_5_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARQOS <= twiddle_h_rsc_0_5_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARPROT <= twiddle_h_rsc_0_5_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARCACHE <= twiddle_h_rsc_0_5_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARBURST <= twiddle_h_rsc_0_5_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARSIZE <= twiddle_h_rsc_0_5_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARLEN <= twiddle_h_rsc_0_5_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_ARADDR <= twiddle_h_rsc_0_5_ARADDR;
  twiddle_h_rsc_0_5_BRESP <= peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_WSTRB <= twiddle_h_rsc_0_5_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_WDATA <= twiddle_h_rsc_0_5_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWREGION <= twiddle_h_rsc_0_5_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWQOS <= twiddle_h_rsc_0_5_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWPROT <= twiddle_h_rsc_0_5_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWCACHE <= twiddle_h_rsc_0_5_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWBURST <= twiddle_h_rsc_0_5_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWSIZE <= twiddle_h_rsc_0_5_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWLEN <= twiddle_h_rsc_0_5_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_AWADDR <= twiddle_h_rsc_0_5_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_5_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_5_i_inst_twiddle_h_rsc_0_5_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_6_i_inst : peaseNTT_core_twiddle_h_rsc_0_6_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_6_s_tdone => twiddle_h_rsc_0_6_s_tdone,
      twiddle_h_rsc_0_6_tr_write_done => twiddle_h_rsc_0_6_tr_write_done,
      twiddle_h_rsc_0_6_RREADY => twiddle_h_rsc_0_6_RREADY,
      twiddle_h_rsc_0_6_RVALID => twiddle_h_rsc_0_6_RVALID,
      twiddle_h_rsc_0_6_RUSER => twiddle_h_rsc_0_6_RUSER,
      twiddle_h_rsc_0_6_RLAST => twiddle_h_rsc_0_6_RLAST,
      twiddle_h_rsc_0_6_RRESP => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_RRESP,
      twiddle_h_rsc_0_6_RDATA => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_RDATA,
      twiddle_h_rsc_0_6_RID => twiddle_h_rsc_0_6_RID,
      twiddle_h_rsc_0_6_ARREADY => twiddle_h_rsc_0_6_ARREADY,
      twiddle_h_rsc_0_6_ARVALID => twiddle_h_rsc_0_6_ARVALID,
      twiddle_h_rsc_0_6_ARUSER => twiddle_h_rsc_0_6_ARUSER,
      twiddle_h_rsc_0_6_ARREGION => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARREGION,
      twiddle_h_rsc_0_6_ARQOS => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARQOS,
      twiddle_h_rsc_0_6_ARPROT => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARPROT,
      twiddle_h_rsc_0_6_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARCACHE,
      twiddle_h_rsc_0_6_ARLOCK => twiddle_h_rsc_0_6_ARLOCK,
      twiddle_h_rsc_0_6_ARBURST => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARBURST,
      twiddle_h_rsc_0_6_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARSIZE,
      twiddle_h_rsc_0_6_ARLEN => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARLEN,
      twiddle_h_rsc_0_6_ARADDR => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARADDR,
      twiddle_h_rsc_0_6_ARID => twiddle_h_rsc_0_6_ARID,
      twiddle_h_rsc_0_6_BREADY => twiddle_h_rsc_0_6_BREADY,
      twiddle_h_rsc_0_6_BVALID => twiddle_h_rsc_0_6_BVALID,
      twiddle_h_rsc_0_6_BUSER => twiddle_h_rsc_0_6_BUSER,
      twiddle_h_rsc_0_6_BRESP => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_BRESP,
      twiddle_h_rsc_0_6_BID => twiddle_h_rsc_0_6_BID,
      twiddle_h_rsc_0_6_WREADY => twiddle_h_rsc_0_6_WREADY,
      twiddle_h_rsc_0_6_WVALID => twiddle_h_rsc_0_6_WVALID,
      twiddle_h_rsc_0_6_WUSER => twiddle_h_rsc_0_6_WUSER,
      twiddle_h_rsc_0_6_WLAST => twiddle_h_rsc_0_6_WLAST,
      twiddle_h_rsc_0_6_WSTRB => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_WSTRB,
      twiddle_h_rsc_0_6_WDATA => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_WDATA,
      twiddle_h_rsc_0_6_AWREADY => twiddle_h_rsc_0_6_AWREADY,
      twiddle_h_rsc_0_6_AWVALID => twiddle_h_rsc_0_6_AWVALID,
      twiddle_h_rsc_0_6_AWUSER => twiddle_h_rsc_0_6_AWUSER,
      twiddle_h_rsc_0_6_AWREGION => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWREGION,
      twiddle_h_rsc_0_6_AWQOS => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWQOS,
      twiddle_h_rsc_0_6_AWPROT => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWPROT,
      twiddle_h_rsc_0_6_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWCACHE,
      twiddle_h_rsc_0_6_AWLOCK => twiddle_h_rsc_0_6_AWLOCK,
      twiddle_h_rsc_0_6_AWBURST => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWBURST,
      twiddle_h_rsc_0_6_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWSIZE,
      twiddle_h_rsc_0_6_AWLEN => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWLEN,
      twiddle_h_rsc_0_6_AWADDR => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWADDR,
      twiddle_h_rsc_0_6_AWID => twiddle_h_rsc_0_6_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_6_i_oswt => reg_twiddle_rsc_0_6_i_oswt_cse,
      twiddle_h_rsc_0_6_i_wen_comp => twiddle_h_rsc_0_6_i_wen_comp,
      twiddle_h_rsc_0_6_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_i_s_raddr_core,
      twiddle_h_rsc_0_6_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_i_s_din_mxwt
    );
  twiddle_h_rsc_0_6_RRESP <= peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_RRESP;
  twiddle_h_rsc_0_6_RDATA <= peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARREGION <= twiddle_h_rsc_0_6_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARQOS <= twiddle_h_rsc_0_6_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARPROT <= twiddle_h_rsc_0_6_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARCACHE <= twiddle_h_rsc_0_6_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARBURST <= twiddle_h_rsc_0_6_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARSIZE <= twiddle_h_rsc_0_6_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARLEN <= twiddle_h_rsc_0_6_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_ARADDR <= twiddle_h_rsc_0_6_ARADDR;
  twiddle_h_rsc_0_6_BRESP <= peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_WSTRB <= twiddle_h_rsc_0_6_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_WDATA <= twiddle_h_rsc_0_6_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWREGION <= twiddle_h_rsc_0_6_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWQOS <= twiddle_h_rsc_0_6_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWPROT <= twiddle_h_rsc_0_6_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWCACHE <= twiddle_h_rsc_0_6_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWBURST <= twiddle_h_rsc_0_6_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWSIZE <= twiddle_h_rsc_0_6_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWLEN <= twiddle_h_rsc_0_6_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_AWADDR <= twiddle_h_rsc_0_6_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_6_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_6_i_inst_twiddle_h_rsc_0_6_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_7_i_inst : peaseNTT_core_twiddle_h_rsc_0_7_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_7_s_tdone => twiddle_h_rsc_0_7_s_tdone,
      twiddle_h_rsc_0_7_tr_write_done => twiddle_h_rsc_0_7_tr_write_done,
      twiddle_h_rsc_0_7_RREADY => twiddle_h_rsc_0_7_RREADY,
      twiddle_h_rsc_0_7_RVALID => twiddle_h_rsc_0_7_RVALID,
      twiddle_h_rsc_0_7_RUSER => twiddle_h_rsc_0_7_RUSER,
      twiddle_h_rsc_0_7_RLAST => twiddle_h_rsc_0_7_RLAST,
      twiddle_h_rsc_0_7_RRESP => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_RRESP,
      twiddle_h_rsc_0_7_RDATA => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_RDATA,
      twiddle_h_rsc_0_7_RID => twiddle_h_rsc_0_7_RID,
      twiddle_h_rsc_0_7_ARREADY => twiddle_h_rsc_0_7_ARREADY,
      twiddle_h_rsc_0_7_ARVALID => twiddle_h_rsc_0_7_ARVALID,
      twiddle_h_rsc_0_7_ARUSER => twiddle_h_rsc_0_7_ARUSER,
      twiddle_h_rsc_0_7_ARREGION => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARREGION,
      twiddle_h_rsc_0_7_ARQOS => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARQOS,
      twiddle_h_rsc_0_7_ARPROT => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARPROT,
      twiddle_h_rsc_0_7_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARCACHE,
      twiddle_h_rsc_0_7_ARLOCK => twiddle_h_rsc_0_7_ARLOCK,
      twiddle_h_rsc_0_7_ARBURST => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARBURST,
      twiddle_h_rsc_0_7_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARSIZE,
      twiddle_h_rsc_0_7_ARLEN => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARLEN,
      twiddle_h_rsc_0_7_ARADDR => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARADDR,
      twiddle_h_rsc_0_7_ARID => twiddle_h_rsc_0_7_ARID,
      twiddle_h_rsc_0_7_BREADY => twiddle_h_rsc_0_7_BREADY,
      twiddle_h_rsc_0_7_BVALID => twiddle_h_rsc_0_7_BVALID,
      twiddle_h_rsc_0_7_BUSER => twiddle_h_rsc_0_7_BUSER,
      twiddle_h_rsc_0_7_BRESP => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_BRESP,
      twiddle_h_rsc_0_7_BID => twiddle_h_rsc_0_7_BID,
      twiddle_h_rsc_0_7_WREADY => twiddle_h_rsc_0_7_WREADY,
      twiddle_h_rsc_0_7_WVALID => twiddle_h_rsc_0_7_WVALID,
      twiddle_h_rsc_0_7_WUSER => twiddle_h_rsc_0_7_WUSER,
      twiddle_h_rsc_0_7_WLAST => twiddle_h_rsc_0_7_WLAST,
      twiddle_h_rsc_0_7_WSTRB => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_WSTRB,
      twiddle_h_rsc_0_7_WDATA => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_WDATA,
      twiddle_h_rsc_0_7_AWREADY => twiddle_h_rsc_0_7_AWREADY,
      twiddle_h_rsc_0_7_AWVALID => twiddle_h_rsc_0_7_AWVALID,
      twiddle_h_rsc_0_7_AWUSER => twiddle_h_rsc_0_7_AWUSER,
      twiddle_h_rsc_0_7_AWREGION => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWREGION,
      twiddle_h_rsc_0_7_AWQOS => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWQOS,
      twiddle_h_rsc_0_7_AWPROT => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWPROT,
      twiddle_h_rsc_0_7_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWCACHE,
      twiddle_h_rsc_0_7_AWLOCK => twiddle_h_rsc_0_7_AWLOCK,
      twiddle_h_rsc_0_7_AWBURST => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWBURST,
      twiddle_h_rsc_0_7_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWSIZE,
      twiddle_h_rsc_0_7_AWLEN => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWLEN,
      twiddle_h_rsc_0_7_AWADDR => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWADDR,
      twiddle_h_rsc_0_7_AWID => twiddle_h_rsc_0_7_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_7_i_oswt => reg_twiddle_rsc_0_7_i_oswt_cse,
      twiddle_h_rsc_0_7_i_wen_comp => twiddle_h_rsc_0_7_i_wen_comp,
      twiddle_h_rsc_0_7_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_i_s_raddr_core,
      twiddle_h_rsc_0_7_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_i_s_din_mxwt
    );
  twiddle_h_rsc_0_7_RRESP <= peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_RRESP;
  twiddle_h_rsc_0_7_RDATA <= peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARREGION <= twiddle_h_rsc_0_7_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARQOS <= twiddle_h_rsc_0_7_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARPROT <= twiddle_h_rsc_0_7_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARCACHE <= twiddle_h_rsc_0_7_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARBURST <= twiddle_h_rsc_0_7_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARSIZE <= twiddle_h_rsc_0_7_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARLEN <= twiddle_h_rsc_0_7_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_ARADDR <= twiddle_h_rsc_0_7_ARADDR;
  twiddle_h_rsc_0_7_BRESP <= peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_WSTRB <= twiddle_h_rsc_0_7_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_WDATA <= twiddle_h_rsc_0_7_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWREGION <= twiddle_h_rsc_0_7_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWQOS <= twiddle_h_rsc_0_7_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWPROT <= twiddle_h_rsc_0_7_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWCACHE <= twiddle_h_rsc_0_7_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWBURST <= twiddle_h_rsc_0_7_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWSIZE <= twiddle_h_rsc_0_7_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWLEN <= twiddle_h_rsc_0_7_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_AWADDR <= twiddle_h_rsc_0_7_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_7_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_7_i_inst_twiddle_h_rsc_0_7_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_8_i_inst : peaseNTT_core_twiddle_h_rsc_0_8_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_8_s_tdone => twiddle_h_rsc_0_8_s_tdone,
      twiddle_h_rsc_0_8_tr_write_done => twiddle_h_rsc_0_8_tr_write_done,
      twiddle_h_rsc_0_8_RREADY => twiddle_h_rsc_0_8_RREADY,
      twiddle_h_rsc_0_8_RVALID => twiddle_h_rsc_0_8_RVALID,
      twiddle_h_rsc_0_8_RUSER => twiddle_h_rsc_0_8_RUSER,
      twiddle_h_rsc_0_8_RLAST => twiddle_h_rsc_0_8_RLAST,
      twiddle_h_rsc_0_8_RRESP => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_RRESP,
      twiddle_h_rsc_0_8_RDATA => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_RDATA,
      twiddle_h_rsc_0_8_RID => twiddle_h_rsc_0_8_RID,
      twiddle_h_rsc_0_8_ARREADY => twiddle_h_rsc_0_8_ARREADY,
      twiddle_h_rsc_0_8_ARVALID => twiddle_h_rsc_0_8_ARVALID,
      twiddle_h_rsc_0_8_ARUSER => twiddle_h_rsc_0_8_ARUSER,
      twiddle_h_rsc_0_8_ARREGION => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARREGION,
      twiddle_h_rsc_0_8_ARQOS => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARQOS,
      twiddle_h_rsc_0_8_ARPROT => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARPROT,
      twiddle_h_rsc_0_8_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARCACHE,
      twiddle_h_rsc_0_8_ARLOCK => twiddle_h_rsc_0_8_ARLOCK,
      twiddle_h_rsc_0_8_ARBURST => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARBURST,
      twiddle_h_rsc_0_8_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARSIZE,
      twiddle_h_rsc_0_8_ARLEN => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARLEN,
      twiddle_h_rsc_0_8_ARADDR => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARADDR,
      twiddle_h_rsc_0_8_ARID => twiddle_h_rsc_0_8_ARID,
      twiddle_h_rsc_0_8_BREADY => twiddle_h_rsc_0_8_BREADY,
      twiddle_h_rsc_0_8_BVALID => twiddle_h_rsc_0_8_BVALID,
      twiddle_h_rsc_0_8_BUSER => twiddle_h_rsc_0_8_BUSER,
      twiddle_h_rsc_0_8_BRESP => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_BRESP,
      twiddle_h_rsc_0_8_BID => twiddle_h_rsc_0_8_BID,
      twiddle_h_rsc_0_8_WREADY => twiddle_h_rsc_0_8_WREADY,
      twiddle_h_rsc_0_8_WVALID => twiddle_h_rsc_0_8_WVALID,
      twiddle_h_rsc_0_8_WUSER => twiddle_h_rsc_0_8_WUSER,
      twiddle_h_rsc_0_8_WLAST => twiddle_h_rsc_0_8_WLAST,
      twiddle_h_rsc_0_8_WSTRB => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_WSTRB,
      twiddle_h_rsc_0_8_WDATA => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_WDATA,
      twiddle_h_rsc_0_8_AWREADY => twiddle_h_rsc_0_8_AWREADY,
      twiddle_h_rsc_0_8_AWVALID => twiddle_h_rsc_0_8_AWVALID,
      twiddle_h_rsc_0_8_AWUSER => twiddle_h_rsc_0_8_AWUSER,
      twiddle_h_rsc_0_8_AWREGION => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWREGION,
      twiddle_h_rsc_0_8_AWQOS => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWQOS,
      twiddle_h_rsc_0_8_AWPROT => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWPROT,
      twiddle_h_rsc_0_8_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWCACHE,
      twiddle_h_rsc_0_8_AWLOCK => twiddle_h_rsc_0_8_AWLOCK,
      twiddle_h_rsc_0_8_AWBURST => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWBURST,
      twiddle_h_rsc_0_8_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWSIZE,
      twiddle_h_rsc_0_8_AWLEN => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWLEN,
      twiddle_h_rsc_0_8_AWADDR => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWADDR,
      twiddle_h_rsc_0_8_AWID => twiddle_h_rsc_0_8_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_8_i_oswt => reg_twiddle_rsc_0_8_i_oswt_cse,
      twiddle_h_rsc_0_8_i_wen_comp => twiddle_h_rsc_0_8_i_wen_comp,
      twiddle_h_rsc_0_8_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_i_s_raddr_core,
      twiddle_h_rsc_0_8_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_i_s_din_mxwt
    );
  twiddle_h_rsc_0_8_RRESP <= peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_RRESP;
  twiddle_h_rsc_0_8_RDATA <= peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARREGION <= twiddle_h_rsc_0_8_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARQOS <= twiddle_h_rsc_0_8_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARPROT <= twiddle_h_rsc_0_8_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARCACHE <= twiddle_h_rsc_0_8_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARBURST <= twiddle_h_rsc_0_8_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARSIZE <= twiddle_h_rsc_0_8_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARLEN <= twiddle_h_rsc_0_8_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_ARADDR <= twiddle_h_rsc_0_8_ARADDR;
  twiddle_h_rsc_0_8_BRESP <= peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_WSTRB <= twiddle_h_rsc_0_8_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_WDATA <= twiddle_h_rsc_0_8_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWREGION <= twiddle_h_rsc_0_8_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWQOS <= twiddle_h_rsc_0_8_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWPROT <= twiddle_h_rsc_0_8_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWCACHE <= twiddle_h_rsc_0_8_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWBURST <= twiddle_h_rsc_0_8_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWSIZE <= twiddle_h_rsc_0_8_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWLEN <= twiddle_h_rsc_0_8_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_AWADDR <= twiddle_h_rsc_0_8_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_8_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_8_i_inst_twiddle_h_rsc_0_8_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_9_i_inst : peaseNTT_core_twiddle_h_rsc_0_9_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_9_s_tdone => twiddle_h_rsc_0_9_s_tdone,
      twiddle_h_rsc_0_9_tr_write_done => twiddle_h_rsc_0_9_tr_write_done,
      twiddle_h_rsc_0_9_RREADY => twiddle_h_rsc_0_9_RREADY,
      twiddle_h_rsc_0_9_RVALID => twiddle_h_rsc_0_9_RVALID,
      twiddle_h_rsc_0_9_RUSER => twiddle_h_rsc_0_9_RUSER,
      twiddle_h_rsc_0_9_RLAST => twiddle_h_rsc_0_9_RLAST,
      twiddle_h_rsc_0_9_RRESP => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_RRESP,
      twiddle_h_rsc_0_9_RDATA => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_RDATA,
      twiddle_h_rsc_0_9_RID => twiddle_h_rsc_0_9_RID,
      twiddle_h_rsc_0_9_ARREADY => twiddle_h_rsc_0_9_ARREADY,
      twiddle_h_rsc_0_9_ARVALID => twiddle_h_rsc_0_9_ARVALID,
      twiddle_h_rsc_0_9_ARUSER => twiddle_h_rsc_0_9_ARUSER,
      twiddle_h_rsc_0_9_ARREGION => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARREGION,
      twiddle_h_rsc_0_9_ARQOS => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARQOS,
      twiddle_h_rsc_0_9_ARPROT => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARPROT,
      twiddle_h_rsc_0_9_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARCACHE,
      twiddle_h_rsc_0_9_ARLOCK => twiddle_h_rsc_0_9_ARLOCK,
      twiddle_h_rsc_0_9_ARBURST => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARBURST,
      twiddle_h_rsc_0_9_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARSIZE,
      twiddle_h_rsc_0_9_ARLEN => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARLEN,
      twiddle_h_rsc_0_9_ARADDR => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARADDR,
      twiddle_h_rsc_0_9_ARID => twiddle_h_rsc_0_9_ARID,
      twiddle_h_rsc_0_9_BREADY => twiddle_h_rsc_0_9_BREADY,
      twiddle_h_rsc_0_9_BVALID => twiddle_h_rsc_0_9_BVALID,
      twiddle_h_rsc_0_9_BUSER => twiddle_h_rsc_0_9_BUSER,
      twiddle_h_rsc_0_9_BRESP => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_BRESP,
      twiddle_h_rsc_0_9_BID => twiddle_h_rsc_0_9_BID,
      twiddle_h_rsc_0_9_WREADY => twiddle_h_rsc_0_9_WREADY,
      twiddle_h_rsc_0_9_WVALID => twiddle_h_rsc_0_9_WVALID,
      twiddle_h_rsc_0_9_WUSER => twiddle_h_rsc_0_9_WUSER,
      twiddle_h_rsc_0_9_WLAST => twiddle_h_rsc_0_9_WLAST,
      twiddle_h_rsc_0_9_WSTRB => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_WSTRB,
      twiddle_h_rsc_0_9_WDATA => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_WDATA,
      twiddle_h_rsc_0_9_AWREADY => twiddle_h_rsc_0_9_AWREADY,
      twiddle_h_rsc_0_9_AWVALID => twiddle_h_rsc_0_9_AWVALID,
      twiddle_h_rsc_0_9_AWUSER => twiddle_h_rsc_0_9_AWUSER,
      twiddle_h_rsc_0_9_AWREGION => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWREGION,
      twiddle_h_rsc_0_9_AWQOS => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWQOS,
      twiddle_h_rsc_0_9_AWPROT => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWPROT,
      twiddle_h_rsc_0_9_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWCACHE,
      twiddle_h_rsc_0_9_AWLOCK => twiddle_h_rsc_0_9_AWLOCK,
      twiddle_h_rsc_0_9_AWBURST => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWBURST,
      twiddle_h_rsc_0_9_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWSIZE,
      twiddle_h_rsc_0_9_AWLEN => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWLEN,
      twiddle_h_rsc_0_9_AWADDR => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWADDR,
      twiddle_h_rsc_0_9_AWID => twiddle_h_rsc_0_9_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_9_i_oswt => reg_twiddle_rsc_0_1_i_oswt_cse,
      twiddle_h_rsc_0_9_i_wen_comp => twiddle_h_rsc_0_9_i_wen_comp,
      twiddle_h_rsc_0_9_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_i_s_raddr_core,
      twiddle_h_rsc_0_9_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_i_s_din_mxwt
    );
  twiddle_h_rsc_0_9_RRESP <= peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_RRESP;
  twiddle_h_rsc_0_9_RDATA <= peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARREGION <= twiddle_h_rsc_0_9_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARQOS <= twiddle_h_rsc_0_9_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARPROT <= twiddle_h_rsc_0_9_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARCACHE <= twiddle_h_rsc_0_9_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARBURST <= twiddle_h_rsc_0_9_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARSIZE <= twiddle_h_rsc_0_9_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARLEN <= twiddle_h_rsc_0_9_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_ARADDR <= twiddle_h_rsc_0_9_ARADDR;
  twiddle_h_rsc_0_9_BRESP <= peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_WSTRB <= twiddle_h_rsc_0_9_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_WDATA <= twiddle_h_rsc_0_9_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWREGION <= twiddle_h_rsc_0_9_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWQOS <= twiddle_h_rsc_0_9_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWPROT <= twiddle_h_rsc_0_9_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWCACHE <= twiddle_h_rsc_0_9_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWBURST <= twiddle_h_rsc_0_9_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWSIZE <= twiddle_h_rsc_0_9_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWLEN <= twiddle_h_rsc_0_9_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_AWADDR <= twiddle_h_rsc_0_9_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_9_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_9_i_inst_twiddle_h_rsc_0_9_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_10_i_inst : peaseNTT_core_twiddle_h_rsc_0_10_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_10_s_tdone => twiddle_h_rsc_0_10_s_tdone,
      twiddle_h_rsc_0_10_tr_write_done => twiddle_h_rsc_0_10_tr_write_done,
      twiddle_h_rsc_0_10_RREADY => twiddle_h_rsc_0_10_RREADY,
      twiddle_h_rsc_0_10_RVALID => twiddle_h_rsc_0_10_RVALID,
      twiddle_h_rsc_0_10_RUSER => twiddle_h_rsc_0_10_RUSER,
      twiddle_h_rsc_0_10_RLAST => twiddle_h_rsc_0_10_RLAST,
      twiddle_h_rsc_0_10_RRESP => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_RRESP,
      twiddle_h_rsc_0_10_RDATA => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_RDATA,
      twiddle_h_rsc_0_10_RID => twiddle_h_rsc_0_10_RID,
      twiddle_h_rsc_0_10_ARREADY => twiddle_h_rsc_0_10_ARREADY,
      twiddle_h_rsc_0_10_ARVALID => twiddle_h_rsc_0_10_ARVALID,
      twiddle_h_rsc_0_10_ARUSER => twiddle_h_rsc_0_10_ARUSER,
      twiddle_h_rsc_0_10_ARREGION => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARREGION,
      twiddle_h_rsc_0_10_ARQOS => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARQOS,
      twiddle_h_rsc_0_10_ARPROT => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARPROT,
      twiddle_h_rsc_0_10_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARCACHE,
      twiddle_h_rsc_0_10_ARLOCK => twiddle_h_rsc_0_10_ARLOCK,
      twiddle_h_rsc_0_10_ARBURST => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARBURST,
      twiddle_h_rsc_0_10_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARSIZE,
      twiddle_h_rsc_0_10_ARLEN => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARLEN,
      twiddle_h_rsc_0_10_ARADDR => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARADDR,
      twiddle_h_rsc_0_10_ARID => twiddle_h_rsc_0_10_ARID,
      twiddle_h_rsc_0_10_BREADY => twiddle_h_rsc_0_10_BREADY,
      twiddle_h_rsc_0_10_BVALID => twiddle_h_rsc_0_10_BVALID,
      twiddle_h_rsc_0_10_BUSER => twiddle_h_rsc_0_10_BUSER,
      twiddle_h_rsc_0_10_BRESP => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_BRESP,
      twiddle_h_rsc_0_10_BID => twiddle_h_rsc_0_10_BID,
      twiddle_h_rsc_0_10_WREADY => twiddle_h_rsc_0_10_WREADY,
      twiddle_h_rsc_0_10_WVALID => twiddle_h_rsc_0_10_WVALID,
      twiddle_h_rsc_0_10_WUSER => twiddle_h_rsc_0_10_WUSER,
      twiddle_h_rsc_0_10_WLAST => twiddle_h_rsc_0_10_WLAST,
      twiddle_h_rsc_0_10_WSTRB => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_WSTRB,
      twiddle_h_rsc_0_10_WDATA => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_WDATA,
      twiddle_h_rsc_0_10_AWREADY => twiddle_h_rsc_0_10_AWREADY,
      twiddle_h_rsc_0_10_AWVALID => twiddle_h_rsc_0_10_AWVALID,
      twiddle_h_rsc_0_10_AWUSER => twiddle_h_rsc_0_10_AWUSER,
      twiddle_h_rsc_0_10_AWREGION => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWREGION,
      twiddle_h_rsc_0_10_AWQOS => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWQOS,
      twiddle_h_rsc_0_10_AWPROT => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWPROT,
      twiddle_h_rsc_0_10_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWCACHE,
      twiddle_h_rsc_0_10_AWLOCK => twiddle_h_rsc_0_10_AWLOCK,
      twiddle_h_rsc_0_10_AWBURST => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWBURST,
      twiddle_h_rsc_0_10_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWSIZE,
      twiddle_h_rsc_0_10_AWLEN => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWLEN,
      twiddle_h_rsc_0_10_AWADDR => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWADDR,
      twiddle_h_rsc_0_10_AWID => twiddle_h_rsc_0_10_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_10_i_oswt => reg_twiddle_rsc_0_2_i_oswt_cse,
      twiddle_h_rsc_0_10_i_wen_comp => twiddle_h_rsc_0_10_i_wen_comp,
      twiddle_h_rsc_0_10_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_i_s_raddr_core,
      twiddle_h_rsc_0_10_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_i_s_din_mxwt
    );
  twiddle_h_rsc_0_10_RRESP <= peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_RRESP;
  twiddle_h_rsc_0_10_RDATA <= peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARREGION <= twiddle_h_rsc_0_10_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARQOS <= twiddle_h_rsc_0_10_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARPROT <= twiddle_h_rsc_0_10_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARCACHE <= twiddle_h_rsc_0_10_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARBURST <= twiddle_h_rsc_0_10_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARSIZE <= twiddle_h_rsc_0_10_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARLEN <= twiddle_h_rsc_0_10_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_ARADDR <= twiddle_h_rsc_0_10_ARADDR;
  twiddle_h_rsc_0_10_BRESP <= peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_WSTRB <= twiddle_h_rsc_0_10_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_WDATA <= twiddle_h_rsc_0_10_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWREGION <= twiddle_h_rsc_0_10_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWQOS <= twiddle_h_rsc_0_10_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWPROT <= twiddle_h_rsc_0_10_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWCACHE <= twiddle_h_rsc_0_10_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWBURST <= twiddle_h_rsc_0_10_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWSIZE <= twiddle_h_rsc_0_10_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWLEN <= twiddle_h_rsc_0_10_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_AWADDR <= twiddle_h_rsc_0_10_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_10_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_10_i_inst_twiddle_h_rsc_0_10_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_11_i_inst : peaseNTT_core_twiddle_h_rsc_0_11_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_11_s_tdone => twiddle_h_rsc_0_11_s_tdone,
      twiddle_h_rsc_0_11_tr_write_done => twiddle_h_rsc_0_11_tr_write_done,
      twiddle_h_rsc_0_11_RREADY => twiddle_h_rsc_0_11_RREADY,
      twiddle_h_rsc_0_11_RVALID => twiddle_h_rsc_0_11_RVALID,
      twiddle_h_rsc_0_11_RUSER => twiddle_h_rsc_0_11_RUSER,
      twiddle_h_rsc_0_11_RLAST => twiddle_h_rsc_0_11_RLAST,
      twiddle_h_rsc_0_11_RRESP => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_RRESP,
      twiddle_h_rsc_0_11_RDATA => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_RDATA,
      twiddle_h_rsc_0_11_RID => twiddle_h_rsc_0_11_RID,
      twiddle_h_rsc_0_11_ARREADY => twiddle_h_rsc_0_11_ARREADY,
      twiddle_h_rsc_0_11_ARVALID => twiddle_h_rsc_0_11_ARVALID,
      twiddle_h_rsc_0_11_ARUSER => twiddle_h_rsc_0_11_ARUSER,
      twiddle_h_rsc_0_11_ARREGION => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARREGION,
      twiddle_h_rsc_0_11_ARQOS => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARQOS,
      twiddle_h_rsc_0_11_ARPROT => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARPROT,
      twiddle_h_rsc_0_11_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARCACHE,
      twiddle_h_rsc_0_11_ARLOCK => twiddle_h_rsc_0_11_ARLOCK,
      twiddle_h_rsc_0_11_ARBURST => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARBURST,
      twiddle_h_rsc_0_11_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARSIZE,
      twiddle_h_rsc_0_11_ARLEN => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARLEN,
      twiddle_h_rsc_0_11_ARADDR => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARADDR,
      twiddle_h_rsc_0_11_ARID => twiddle_h_rsc_0_11_ARID,
      twiddle_h_rsc_0_11_BREADY => twiddle_h_rsc_0_11_BREADY,
      twiddle_h_rsc_0_11_BVALID => twiddle_h_rsc_0_11_BVALID,
      twiddle_h_rsc_0_11_BUSER => twiddle_h_rsc_0_11_BUSER,
      twiddle_h_rsc_0_11_BRESP => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_BRESP,
      twiddle_h_rsc_0_11_BID => twiddle_h_rsc_0_11_BID,
      twiddle_h_rsc_0_11_WREADY => twiddle_h_rsc_0_11_WREADY,
      twiddle_h_rsc_0_11_WVALID => twiddle_h_rsc_0_11_WVALID,
      twiddle_h_rsc_0_11_WUSER => twiddle_h_rsc_0_11_WUSER,
      twiddle_h_rsc_0_11_WLAST => twiddle_h_rsc_0_11_WLAST,
      twiddle_h_rsc_0_11_WSTRB => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_WSTRB,
      twiddle_h_rsc_0_11_WDATA => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_WDATA,
      twiddle_h_rsc_0_11_AWREADY => twiddle_h_rsc_0_11_AWREADY,
      twiddle_h_rsc_0_11_AWVALID => twiddle_h_rsc_0_11_AWVALID,
      twiddle_h_rsc_0_11_AWUSER => twiddle_h_rsc_0_11_AWUSER,
      twiddle_h_rsc_0_11_AWREGION => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWREGION,
      twiddle_h_rsc_0_11_AWQOS => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWQOS,
      twiddle_h_rsc_0_11_AWPROT => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWPROT,
      twiddle_h_rsc_0_11_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWCACHE,
      twiddle_h_rsc_0_11_AWLOCK => twiddle_h_rsc_0_11_AWLOCK,
      twiddle_h_rsc_0_11_AWBURST => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWBURST,
      twiddle_h_rsc_0_11_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWSIZE,
      twiddle_h_rsc_0_11_AWLEN => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWLEN,
      twiddle_h_rsc_0_11_AWADDR => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWADDR,
      twiddle_h_rsc_0_11_AWID => twiddle_h_rsc_0_11_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_11_i_oswt => reg_twiddle_rsc_0_3_i_oswt_cse,
      twiddle_h_rsc_0_11_i_wen_comp => twiddle_h_rsc_0_11_i_wen_comp,
      twiddle_h_rsc_0_11_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_i_s_raddr_core,
      twiddle_h_rsc_0_11_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_i_s_din_mxwt
    );
  twiddle_h_rsc_0_11_RRESP <= peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_RRESP;
  twiddle_h_rsc_0_11_RDATA <= peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARREGION <= twiddle_h_rsc_0_11_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARQOS <= twiddle_h_rsc_0_11_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARPROT <= twiddle_h_rsc_0_11_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARCACHE <= twiddle_h_rsc_0_11_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARBURST <= twiddle_h_rsc_0_11_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARSIZE <= twiddle_h_rsc_0_11_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARLEN <= twiddle_h_rsc_0_11_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_ARADDR <= twiddle_h_rsc_0_11_ARADDR;
  twiddle_h_rsc_0_11_BRESP <= peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_WSTRB <= twiddle_h_rsc_0_11_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_WDATA <= twiddle_h_rsc_0_11_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWREGION <= twiddle_h_rsc_0_11_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWQOS <= twiddle_h_rsc_0_11_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWPROT <= twiddle_h_rsc_0_11_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWCACHE <= twiddle_h_rsc_0_11_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWBURST <= twiddle_h_rsc_0_11_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWSIZE <= twiddle_h_rsc_0_11_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWLEN <= twiddle_h_rsc_0_11_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_AWADDR <= twiddle_h_rsc_0_11_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_11_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_11_i_inst_twiddle_h_rsc_0_11_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_12_i_inst : peaseNTT_core_twiddle_h_rsc_0_12_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_12_s_tdone => twiddle_h_rsc_0_12_s_tdone,
      twiddle_h_rsc_0_12_tr_write_done => twiddle_h_rsc_0_12_tr_write_done,
      twiddle_h_rsc_0_12_RREADY => twiddle_h_rsc_0_12_RREADY,
      twiddle_h_rsc_0_12_RVALID => twiddle_h_rsc_0_12_RVALID,
      twiddle_h_rsc_0_12_RUSER => twiddle_h_rsc_0_12_RUSER,
      twiddle_h_rsc_0_12_RLAST => twiddle_h_rsc_0_12_RLAST,
      twiddle_h_rsc_0_12_RRESP => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_RRESP,
      twiddle_h_rsc_0_12_RDATA => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_RDATA,
      twiddle_h_rsc_0_12_RID => twiddle_h_rsc_0_12_RID,
      twiddle_h_rsc_0_12_ARREADY => twiddle_h_rsc_0_12_ARREADY,
      twiddle_h_rsc_0_12_ARVALID => twiddle_h_rsc_0_12_ARVALID,
      twiddle_h_rsc_0_12_ARUSER => twiddle_h_rsc_0_12_ARUSER,
      twiddle_h_rsc_0_12_ARREGION => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARREGION,
      twiddle_h_rsc_0_12_ARQOS => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARQOS,
      twiddle_h_rsc_0_12_ARPROT => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARPROT,
      twiddle_h_rsc_0_12_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARCACHE,
      twiddle_h_rsc_0_12_ARLOCK => twiddle_h_rsc_0_12_ARLOCK,
      twiddle_h_rsc_0_12_ARBURST => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARBURST,
      twiddle_h_rsc_0_12_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARSIZE,
      twiddle_h_rsc_0_12_ARLEN => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARLEN,
      twiddle_h_rsc_0_12_ARADDR => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARADDR,
      twiddle_h_rsc_0_12_ARID => twiddle_h_rsc_0_12_ARID,
      twiddle_h_rsc_0_12_BREADY => twiddle_h_rsc_0_12_BREADY,
      twiddle_h_rsc_0_12_BVALID => twiddle_h_rsc_0_12_BVALID,
      twiddle_h_rsc_0_12_BUSER => twiddle_h_rsc_0_12_BUSER,
      twiddle_h_rsc_0_12_BRESP => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_BRESP,
      twiddle_h_rsc_0_12_BID => twiddle_h_rsc_0_12_BID,
      twiddle_h_rsc_0_12_WREADY => twiddle_h_rsc_0_12_WREADY,
      twiddle_h_rsc_0_12_WVALID => twiddle_h_rsc_0_12_WVALID,
      twiddle_h_rsc_0_12_WUSER => twiddle_h_rsc_0_12_WUSER,
      twiddle_h_rsc_0_12_WLAST => twiddle_h_rsc_0_12_WLAST,
      twiddle_h_rsc_0_12_WSTRB => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_WSTRB,
      twiddle_h_rsc_0_12_WDATA => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_WDATA,
      twiddle_h_rsc_0_12_AWREADY => twiddle_h_rsc_0_12_AWREADY,
      twiddle_h_rsc_0_12_AWVALID => twiddle_h_rsc_0_12_AWVALID,
      twiddle_h_rsc_0_12_AWUSER => twiddle_h_rsc_0_12_AWUSER,
      twiddle_h_rsc_0_12_AWREGION => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWREGION,
      twiddle_h_rsc_0_12_AWQOS => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWQOS,
      twiddle_h_rsc_0_12_AWPROT => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWPROT,
      twiddle_h_rsc_0_12_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWCACHE,
      twiddle_h_rsc_0_12_AWLOCK => twiddle_h_rsc_0_12_AWLOCK,
      twiddle_h_rsc_0_12_AWBURST => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWBURST,
      twiddle_h_rsc_0_12_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWSIZE,
      twiddle_h_rsc_0_12_AWLEN => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWLEN,
      twiddle_h_rsc_0_12_AWADDR => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWADDR,
      twiddle_h_rsc_0_12_AWID => twiddle_h_rsc_0_12_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_12_i_oswt => reg_twiddle_rsc_0_4_i_oswt_cse,
      twiddle_h_rsc_0_12_i_wen_comp => twiddle_h_rsc_0_12_i_wen_comp,
      twiddle_h_rsc_0_12_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_i_s_raddr_core,
      twiddle_h_rsc_0_12_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_i_s_din_mxwt
    );
  twiddle_h_rsc_0_12_RRESP <= peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_RRESP;
  twiddle_h_rsc_0_12_RDATA <= peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARREGION <= twiddle_h_rsc_0_12_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARQOS <= twiddle_h_rsc_0_12_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARPROT <= twiddle_h_rsc_0_12_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARCACHE <= twiddle_h_rsc_0_12_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARBURST <= twiddle_h_rsc_0_12_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARSIZE <= twiddle_h_rsc_0_12_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARLEN <= twiddle_h_rsc_0_12_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_ARADDR <= twiddle_h_rsc_0_12_ARADDR;
  twiddle_h_rsc_0_12_BRESP <= peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_WSTRB <= twiddle_h_rsc_0_12_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_WDATA <= twiddle_h_rsc_0_12_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWREGION <= twiddle_h_rsc_0_12_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWQOS <= twiddle_h_rsc_0_12_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWPROT <= twiddle_h_rsc_0_12_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWCACHE <= twiddle_h_rsc_0_12_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWBURST <= twiddle_h_rsc_0_12_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWSIZE <= twiddle_h_rsc_0_12_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWLEN <= twiddle_h_rsc_0_12_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_AWADDR <= twiddle_h_rsc_0_12_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_12_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_12_i_inst_twiddle_h_rsc_0_12_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_13_i_inst : peaseNTT_core_twiddle_h_rsc_0_13_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_13_s_tdone => twiddle_h_rsc_0_13_s_tdone,
      twiddle_h_rsc_0_13_tr_write_done => twiddle_h_rsc_0_13_tr_write_done,
      twiddle_h_rsc_0_13_RREADY => twiddle_h_rsc_0_13_RREADY,
      twiddle_h_rsc_0_13_RVALID => twiddle_h_rsc_0_13_RVALID,
      twiddle_h_rsc_0_13_RUSER => twiddle_h_rsc_0_13_RUSER,
      twiddle_h_rsc_0_13_RLAST => twiddle_h_rsc_0_13_RLAST,
      twiddle_h_rsc_0_13_RRESP => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_RRESP,
      twiddle_h_rsc_0_13_RDATA => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_RDATA,
      twiddle_h_rsc_0_13_RID => twiddle_h_rsc_0_13_RID,
      twiddle_h_rsc_0_13_ARREADY => twiddle_h_rsc_0_13_ARREADY,
      twiddle_h_rsc_0_13_ARVALID => twiddle_h_rsc_0_13_ARVALID,
      twiddle_h_rsc_0_13_ARUSER => twiddle_h_rsc_0_13_ARUSER,
      twiddle_h_rsc_0_13_ARREGION => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARREGION,
      twiddle_h_rsc_0_13_ARQOS => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARQOS,
      twiddle_h_rsc_0_13_ARPROT => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARPROT,
      twiddle_h_rsc_0_13_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARCACHE,
      twiddle_h_rsc_0_13_ARLOCK => twiddle_h_rsc_0_13_ARLOCK,
      twiddle_h_rsc_0_13_ARBURST => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARBURST,
      twiddle_h_rsc_0_13_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARSIZE,
      twiddle_h_rsc_0_13_ARLEN => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARLEN,
      twiddle_h_rsc_0_13_ARADDR => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARADDR,
      twiddle_h_rsc_0_13_ARID => twiddle_h_rsc_0_13_ARID,
      twiddle_h_rsc_0_13_BREADY => twiddle_h_rsc_0_13_BREADY,
      twiddle_h_rsc_0_13_BVALID => twiddle_h_rsc_0_13_BVALID,
      twiddle_h_rsc_0_13_BUSER => twiddle_h_rsc_0_13_BUSER,
      twiddle_h_rsc_0_13_BRESP => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_BRESP,
      twiddle_h_rsc_0_13_BID => twiddle_h_rsc_0_13_BID,
      twiddle_h_rsc_0_13_WREADY => twiddle_h_rsc_0_13_WREADY,
      twiddle_h_rsc_0_13_WVALID => twiddle_h_rsc_0_13_WVALID,
      twiddle_h_rsc_0_13_WUSER => twiddle_h_rsc_0_13_WUSER,
      twiddle_h_rsc_0_13_WLAST => twiddle_h_rsc_0_13_WLAST,
      twiddle_h_rsc_0_13_WSTRB => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_WSTRB,
      twiddle_h_rsc_0_13_WDATA => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_WDATA,
      twiddle_h_rsc_0_13_AWREADY => twiddle_h_rsc_0_13_AWREADY,
      twiddle_h_rsc_0_13_AWVALID => twiddle_h_rsc_0_13_AWVALID,
      twiddle_h_rsc_0_13_AWUSER => twiddle_h_rsc_0_13_AWUSER,
      twiddle_h_rsc_0_13_AWREGION => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWREGION,
      twiddle_h_rsc_0_13_AWQOS => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWQOS,
      twiddle_h_rsc_0_13_AWPROT => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWPROT,
      twiddle_h_rsc_0_13_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWCACHE,
      twiddle_h_rsc_0_13_AWLOCK => twiddle_h_rsc_0_13_AWLOCK,
      twiddle_h_rsc_0_13_AWBURST => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWBURST,
      twiddle_h_rsc_0_13_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWSIZE,
      twiddle_h_rsc_0_13_AWLEN => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWLEN,
      twiddle_h_rsc_0_13_AWADDR => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWADDR,
      twiddle_h_rsc_0_13_AWID => twiddle_h_rsc_0_13_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_13_i_oswt => reg_twiddle_rsc_0_5_i_oswt_cse,
      twiddle_h_rsc_0_13_i_wen_comp => twiddle_h_rsc_0_13_i_wen_comp,
      twiddle_h_rsc_0_13_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_i_s_raddr_core,
      twiddle_h_rsc_0_13_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_i_s_din_mxwt
    );
  twiddle_h_rsc_0_13_RRESP <= peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_RRESP;
  twiddle_h_rsc_0_13_RDATA <= peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARREGION <= twiddle_h_rsc_0_13_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARQOS <= twiddle_h_rsc_0_13_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARPROT <= twiddle_h_rsc_0_13_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARCACHE <= twiddle_h_rsc_0_13_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARBURST <= twiddle_h_rsc_0_13_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARSIZE <= twiddle_h_rsc_0_13_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARLEN <= twiddle_h_rsc_0_13_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_ARADDR <= twiddle_h_rsc_0_13_ARADDR;
  twiddle_h_rsc_0_13_BRESP <= peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_WSTRB <= twiddle_h_rsc_0_13_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_WDATA <= twiddle_h_rsc_0_13_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWREGION <= twiddle_h_rsc_0_13_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWQOS <= twiddle_h_rsc_0_13_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWPROT <= twiddle_h_rsc_0_13_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWCACHE <= twiddle_h_rsc_0_13_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWBURST <= twiddle_h_rsc_0_13_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWSIZE <= twiddle_h_rsc_0_13_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWLEN <= twiddle_h_rsc_0_13_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_AWADDR <= twiddle_h_rsc_0_13_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_13_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_13_i_inst_twiddle_h_rsc_0_13_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_14_i_inst : peaseNTT_core_twiddle_h_rsc_0_14_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_14_s_tdone => twiddle_h_rsc_0_14_s_tdone,
      twiddle_h_rsc_0_14_tr_write_done => twiddle_h_rsc_0_14_tr_write_done,
      twiddle_h_rsc_0_14_RREADY => twiddle_h_rsc_0_14_RREADY,
      twiddle_h_rsc_0_14_RVALID => twiddle_h_rsc_0_14_RVALID,
      twiddle_h_rsc_0_14_RUSER => twiddle_h_rsc_0_14_RUSER,
      twiddle_h_rsc_0_14_RLAST => twiddle_h_rsc_0_14_RLAST,
      twiddle_h_rsc_0_14_RRESP => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_RRESP,
      twiddle_h_rsc_0_14_RDATA => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_RDATA,
      twiddle_h_rsc_0_14_RID => twiddle_h_rsc_0_14_RID,
      twiddle_h_rsc_0_14_ARREADY => twiddle_h_rsc_0_14_ARREADY,
      twiddle_h_rsc_0_14_ARVALID => twiddle_h_rsc_0_14_ARVALID,
      twiddle_h_rsc_0_14_ARUSER => twiddle_h_rsc_0_14_ARUSER,
      twiddle_h_rsc_0_14_ARREGION => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARREGION,
      twiddle_h_rsc_0_14_ARQOS => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARQOS,
      twiddle_h_rsc_0_14_ARPROT => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARPROT,
      twiddle_h_rsc_0_14_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARCACHE,
      twiddle_h_rsc_0_14_ARLOCK => twiddle_h_rsc_0_14_ARLOCK,
      twiddle_h_rsc_0_14_ARBURST => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARBURST,
      twiddle_h_rsc_0_14_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARSIZE,
      twiddle_h_rsc_0_14_ARLEN => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARLEN,
      twiddle_h_rsc_0_14_ARADDR => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARADDR,
      twiddle_h_rsc_0_14_ARID => twiddle_h_rsc_0_14_ARID,
      twiddle_h_rsc_0_14_BREADY => twiddle_h_rsc_0_14_BREADY,
      twiddle_h_rsc_0_14_BVALID => twiddle_h_rsc_0_14_BVALID,
      twiddle_h_rsc_0_14_BUSER => twiddle_h_rsc_0_14_BUSER,
      twiddle_h_rsc_0_14_BRESP => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_BRESP,
      twiddle_h_rsc_0_14_BID => twiddle_h_rsc_0_14_BID,
      twiddle_h_rsc_0_14_WREADY => twiddle_h_rsc_0_14_WREADY,
      twiddle_h_rsc_0_14_WVALID => twiddle_h_rsc_0_14_WVALID,
      twiddle_h_rsc_0_14_WUSER => twiddle_h_rsc_0_14_WUSER,
      twiddle_h_rsc_0_14_WLAST => twiddle_h_rsc_0_14_WLAST,
      twiddle_h_rsc_0_14_WSTRB => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_WSTRB,
      twiddle_h_rsc_0_14_WDATA => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_WDATA,
      twiddle_h_rsc_0_14_AWREADY => twiddle_h_rsc_0_14_AWREADY,
      twiddle_h_rsc_0_14_AWVALID => twiddle_h_rsc_0_14_AWVALID,
      twiddle_h_rsc_0_14_AWUSER => twiddle_h_rsc_0_14_AWUSER,
      twiddle_h_rsc_0_14_AWREGION => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWREGION,
      twiddle_h_rsc_0_14_AWQOS => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWQOS,
      twiddle_h_rsc_0_14_AWPROT => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWPROT,
      twiddle_h_rsc_0_14_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWCACHE,
      twiddle_h_rsc_0_14_AWLOCK => twiddle_h_rsc_0_14_AWLOCK,
      twiddle_h_rsc_0_14_AWBURST => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWBURST,
      twiddle_h_rsc_0_14_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWSIZE,
      twiddle_h_rsc_0_14_AWLEN => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWLEN,
      twiddle_h_rsc_0_14_AWADDR => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWADDR,
      twiddle_h_rsc_0_14_AWID => twiddle_h_rsc_0_14_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_14_i_oswt => reg_twiddle_rsc_0_6_i_oswt_cse,
      twiddle_h_rsc_0_14_i_wen_comp => twiddle_h_rsc_0_14_i_wen_comp,
      twiddle_h_rsc_0_14_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_i_s_raddr_core,
      twiddle_h_rsc_0_14_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_i_s_din_mxwt
    );
  twiddle_h_rsc_0_14_RRESP <= peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_RRESP;
  twiddle_h_rsc_0_14_RDATA <= peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARREGION <= twiddle_h_rsc_0_14_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARQOS <= twiddle_h_rsc_0_14_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARPROT <= twiddle_h_rsc_0_14_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARCACHE <= twiddle_h_rsc_0_14_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARBURST <= twiddle_h_rsc_0_14_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARSIZE <= twiddle_h_rsc_0_14_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARLEN <= twiddle_h_rsc_0_14_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_ARADDR <= twiddle_h_rsc_0_14_ARADDR;
  twiddle_h_rsc_0_14_BRESP <= peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_WSTRB <= twiddle_h_rsc_0_14_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_WDATA <= twiddle_h_rsc_0_14_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWREGION <= twiddle_h_rsc_0_14_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWQOS <= twiddle_h_rsc_0_14_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWPROT <= twiddle_h_rsc_0_14_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWCACHE <= twiddle_h_rsc_0_14_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWBURST <= twiddle_h_rsc_0_14_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWSIZE <= twiddle_h_rsc_0_14_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWLEN <= twiddle_h_rsc_0_14_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_AWADDR <= twiddle_h_rsc_0_14_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_14_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_14_i_inst_twiddle_h_rsc_0_14_i_s_din_mxwt;

  peaseNTT_core_twiddle_h_rsc_0_15_i_inst : peaseNTT_core_twiddle_h_rsc_0_15_i
    PORT MAP(
      clk => clk,
      rst => rst,
      twiddle_h_rsc_0_15_s_tdone => twiddle_h_rsc_0_15_s_tdone,
      twiddle_h_rsc_0_15_tr_write_done => twiddle_h_rsc_0_15_tr_write_done,
      twiddle_h_rsc_0_15_RREADY => twiddle_h_rsc_0_15_RREADY,
      twiddle_h_rsc_0_15_RVALID => twiddle_h_rsc_0_15_RVALID,
      twiddle_h_rsc_0_15_RUSER => twiddle_h_rsc_0_15_RUSER,
      twiddle_h_rsc_0_15_RLAST => twiddle_h_rsc_0_15_RLAST,
      twiddle_h_rsc_0_15_RRESP => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_RRESP,
      twiddle_h_rsc_0_15_RDATA => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_RDATA,
      twiddle_h_rsc_0_15_RID => twiddle_h_rsc_0_15_RID,
      twiddle_h_rsc_0_15_ARREADY => twiddle_h_rsc_0_15_ARREADY,
      twiddle_h_rsc_0_15_ARVALID => twiddle_h_rsc_0_15_ARVALID,
      twiddle_h_rsc_0_15_ARUSER => twiddle_h_rsc_0_15_ARUSER,
      twiddle_h_rsc_0_15_ARREGION => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARREGION,
      twiddle_h_rsc_0_15_ARQOS => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARQOS,
      twiddle_h_rsc_0_15_ARPROT => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARPROT,
      twiddle_h_rsc_0_15_ARCACHE => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARCACHE,
      twiddle_h_rsc_0_15_ARLOCK => twiddle_h_rsc_0_15_ARLOCK,
      twiddle_h_rsc_0_15_ARBURST => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARBURST,
      twiddle_h_rsc_0_15_ARSIZE => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARSIZE,
      twiddle_h_rsc_0_15_ARLEN => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARLEN,
      twiddle_h_rsc_0_15_ARADDR => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARADDR,
      twiddle_h_rsc_0_15_ARID => twiddle_h_rsc_0_15_ARID,
      twiddle_h_rsc_0_15_BREADY => twiddle_h_rsc_0_15_BREADY,
      twiddle_h_rsc_0_15_BVALID => twiddle_h_rsc_0_15_BVALID,
      twiddle_h_rsc_0_15_BUSER => twiddle_h_rsc_0_15_BUSER,
      twiddle_h_rsc_0_15_BRESP => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_BRESP,
      twiddle_h_rsc_0_15_BID => twiddle_h_rsc_0_15_BID,
      twiddle_h_rsc_0_15_WREADY => twiddle_h_rsc_0_15_WREADY,
      twiddle_h_rsc_0_15_WVALID => twiddle_h_rsc_0_15_WVALID,
      twiddle_h_rsc_0_15_WUSER => twiddle_h_rsc_0_15_WUSER,
      twiddle_h_rsc_0_15_WLAST => twiddle_h_rsc_0_15_WLAST,
      twiddle_h_rsc_0_15_WSTRB => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_WSTRB,
      twiddle_h_rsc_0_15_WDATA => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_WDATA,
      twiddle_h_rsc_0_15_AWREADY => twiddle_h_rsc_0_15_AWREADY,
      twiddle_h_rsc_0_15_AWVALID => twiddle_h_rsc_0_15_AWVALID,
      twiddle_h_rsc_0_15_AWUSER => twiddle_h_rsc_0_15_AWUSER,
      twiddle_h_rsc_0_15_AWREGION => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWREGION,
      twiddle_h_rsc_0_15_AWQOS => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWQOS,
      twiddle_h_rsc_0_15_AWPROT => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWPROT,
      twiddle_h_rsc_0_15_AWCACHE => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWCACHE,
      twiddle_h_rsc_0_15_AWLOCK => twiddle_h_rsc_0_15_AWLOCK,
      twiddle_h_rsc_0_15_AWBURST => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWBURST,
      twiddle_h_rsc_0_15_AWSIZE => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWSIZE,
      twiddle_h_rsc_0_15_AWLEN => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWLEN,
      twiddle_h_rsc_0_15_AWADDR => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWADDR,
      twiddle_h_rsc_0_15_AWID => twiddle_h_rsc_0_15_AWID,
      core_wen => core_wen,
      twiddle_h_rsc_0_15_i_oswt => reg_twiddle_rsc_0_7_i_oswt_cse,
      twiddle_h_rsc_0_15_i_wen_comp => twiddle_h_rsc_0_15_i_wen_comp,
      twiddle_h_rsc_0_15_i_s_raddr_core => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_i_s_raddr_core,
      twiddle_h_rsc_0_15_i_s_din_mxwt => peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_i_s_din_mxwt
    );
  twiddle_h_rsc_0_15_RRESP <= peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_RRESP;
  twiddle_h_rsc_0_15_RDATA <= peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_RDATA;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARREGION <= twiddle_h_rsc_0_15_ARREGION;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARQOS <= twiddle_h_rsc_0_15_ARQOS;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARPROT <= twiddle_h_rsc_0_15_ARPROT;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARCACHE <= twiddle_h_rsc_0_15_ARCACHE;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARBURST <= twiddle_h_rsc_0_15_ARBURST;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARSIZE <= twiddle_h_rsc_0_15_ARSIZE;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARLEN <= twiddle_h_rsc_0_15_ARLEN;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_ARADDR <= twiddle_h_rsc_0_15_ARADDR;
  twiddle_h_rsc_0_15_BRESP <= peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_BRESP;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_WSTRB <= twiddle_h_rsc_0_15_WSTRB;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_WDATA <= twiddle_h_rsc_0_15_WDATA;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWREGION <= twiddle_h_rsc_0_15_AWREGION;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWQOS <= twiddle_h_rsc_0_15_AWQOS;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWPROT <= twiddle_h_rsc_0_15_AWPROT;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWCACHE <= twiddle_h_rsc_0_15_AWCACHE;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWBURST <= twiddle_h_rsc_0_15_AWBURST;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWSIZE <= twiddle_h_rsc_0_15_AWSIZE;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWLEN <= twiddle_h_rsc_0_15_AWLEN;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_AWADDR <= twiddle_h_rsc_0_15_AWADDR;
  peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_i_s_raddr_core <= STD_LOGIC_VECTOR(UNSIGNED'(
      "0") & UNSIGNED(reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse));
  twiddle_h_rsc_0_15_i_s_din_mxwt <= peaseNTT_core_twiddle_h_rsc_0_15_i_inst_twiddle_h_rsc_0_15_i_s_din_mxwt;

  peaseNTT_core_xt_rsc_triosy_1_31_obj_inst : peaseNTT_core_xt_rsc_triosy_1_31_obj
    PORT MAP(
      xt_rsc_triosy_1_31_lz => xt_rsc_triosy_1_31_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_31_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_30_obj_inst : peaseNTT_core_xt_rsc_triosy_1_30_obj
    PORT MAP(
      xt_rsc_triosy_1_30_lz => xt_rsc_triosy_1_30_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_30_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_29_obj_inst : peaseNTT_core_xt_rsc_triosy_1_29_obj
    PORT MAP(
      xt_rsc_triosy_1_29_lz => xt_rsc_triosy_1_29_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_29_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_28_obj_inst : peaseNTT_core_xt_rsc_triosy_1_28_obj
    PORT MAP(
      xt_rsc_triosy_1_28_lz => xt_rsc_triosy_1_28_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_28_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_27_obj_inst : peaseNTT_core_xt_rsc_triosy_1_27_obj
    PORT MAP(
      xt_rsc_triosy_1_27_lz => xt_rsc_triosy_1_27_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_27_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_26_obj_inst : peaseNTT_core_xt_rsc_triosy_1_26_obj
    PORT MAP(
      xt_rsc_triosy_1_26_lz => xt_rsc_triosy_1_26_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_26_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_25_obj_inst : peaseNTT_core_xt_rsc_triosy_1_25_obj
    PORT MAP(
      xt_rsc_triosy_1_25_lz => xt_rsc_triosy_1_25_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_25_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_24_obj_inst : peaseNTT_core_xt_rsc_triosy_1_24_obj
    PORT MAP(
      xt_rsc_triosy_1_24_lz => xt_rsc_triosy_1_24_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_24_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_23_obj_inst : peaseNTT_core_xt_rsc_triosy_1_23_obj
    PORT MAP(
      xt_rsc_triosy_1_23_lz => xt_rsc_triosy_1_23_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_23_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_22_obj_inst : peaseNTT_core_xt_rsc_triosy_1_22_obj
    PORT MAP(
      xt_rsc_triosy_1_22_lz => xt_rsc_triosy_1_22_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_22_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_21_obj_inst : peaseNTT_core_xt_rsc_triosy_1_21_obj
    PORT MAP(
      xt_rsc_triosy_1_21_lz => xt_rsc_triosy_1_21_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_21_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_20_obj_inst : peaseNTT_core_xt_rsc_triosy_1_20_obj
    PORT MAP(
      xt_rsc_triosy_1_20_lz => xt_rsc_triosy_1_20_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_20_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_19_obj_inst : peaseNTT_core_xt_rsc_triosy_1_19_obj
    PORT MAP(
      xt_rsc_triosy_1_19_lz => xt_rsc_triosy_1_19_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_19_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_18_obj_inst : peaseNTT_core_xt_rsc_triosy_1_18_obj
    PORT MAP(
      xt_rsc_triosy_1_18_lz => xt_rsc_triosy_1_18_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_18_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_17_obj_inst : peaseNTT_core_xt_rsc_triosy_1_17_obj
    PORT MAP(
      xt_rsc_triosy_1_17_lz => xt_rsc_triosy_1_17_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_17_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_16_obj_inst : peaseNTT_core_xt_rsc_triosy_1_16_obj
    PORT MAP(
      xt_rsc_triosy_1_16_lz => xt_rsc_triosy_1_16_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_16_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_15_obj_inst : peaseNTT_core_xt_rsc_triosy_1_15_obj
    PORT MAP(
      xt_rsc_triosy_1_15_lz => xt_rsc_triosy_1_15_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_15_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_14_obj_inst : peaseNTT_core_xt_rsc_triosy_1_14_obj
    PORT MAP(
      xt_rsc_triosy_1_14_lz => xt_rsc_triosy_1_14_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_14_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_13_obj_inst : peaseNTT_core_xt_rsc_triosy_1_13_obj
    PORT MAP(
      xt_rsc_triosy_1_13_lz => xt_rsc_triosy_1_13_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_13_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_12_obj_inst : peaseNTT_core_xt_rsc_triosy_1_12_obj
    PORT MAP(
      xt_rsc_triosy_1_12_lz => xt_rsc_triosy_1_12_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_12_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_11_obj_inst : peaseNTT_core_xt_rsc_triosy_1_11_obj
    PORT MAP(
      xt_rsc_triosy_1_11_lz => xt_rsc_triosy_1_11_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_11_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_10_obj_inst : peaseNTT_core_xt_rsc_triosy_1_10_obj
    PORT MAP(
      xt_rsc_triosy_1_10_lz => xt_rsc_triosy_1_10_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_10_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_9_obj_inst : peaseNTT_core_xt_rsc_triosy_1_9_obj
    PORT MAP(
      xt_rsc_triosy_1_9_lz => xt_rsc_triosy_1_9_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_9_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_8_obj_inst : peaseNTT_core_xt_rsc_triosy_1_8_obj
    PORT MAP(
      xt_rsc_triosy_1_8_lz => xt_rsc_triosy_1_8_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_8_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_7_obj_inst : peaseNTT_core_xt_rsc_triosy_1_7_obj
    PORT MAP(
      xt_rsc_triosy_1_7_lz => xt_rsc_triosy_1_7_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_7_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_6_obj_inst : peaseNTT_core_xt_rsc_triosy_1_6_obj
    PORT MAP(
      xt_rsc_triosy_1_6_lz => xt_rsc_triosy_1_6_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_6_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_5_obj_inst : peaseNTT_core_xt_rsc_triosy_1_5_obj
    PORT MAP(
      xt_rsc_triosy_1_5_lz => xt_rsc_triosy_1_5_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_5_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_4_obj_inst : peaseNTT_core_xt_rsc_triosy_1_4_obj
    PORT MAP(
      xt_rsc_triosy_1_4_lz => xt_rsc_triosy_1_4_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_4_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_3_obj_inst : peaseNTT_core_xt_rsc_triosy_1_3_obj
    PORT MAP(
      xt_rsc_triosy_1_3_lz => xt_rsc_triosy_1_3_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_3_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_2_obj_inst : peaseNTT_core_xt_rsc_triosy_1_2_obj
    PORT MAP(
      xt_rsc_triosy_1_2_lz => xt_rsc_triosy_1_2_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_2_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_1_obj_inst : peaseNTT_core_xt_rsc_triosy_1_1_obj
    PORT MAP(
      xt_rsc_triosy_1_1_lz => xt_rsc_triosy_1_1_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_1_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_1_0_obj_inst : peaseNTT_core_xt_rsc_triosy_1_0_obj
    PORT MAP(
      xt_rsc_triosy_1_0_lz => xt_rsc_triosy_1_0_lz,
      core_wten => core_wten,
      xt_rsc_triosy_1_0_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_31_obj_inst : peaseNTT_core_xt_rsc_triosy_0_31_obj
    PORT MAP(
      xt_rsc_triosy_0_31_lz => xt_rsc_triosy_0_31_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_31_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_30_obj_inst : peaseNTT_core_xt_rsc_triosy_0_30_obj
    PORT MAP(
      xt_rsc_triosy_0_30_lz => xt_rsc_triosy_0_30_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_30_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_29_obj_inst : peaseNTT_core_xt_rsc_triosy_0_29_obj
    PORT MAP(
      xt_rsc_triosy_0_29_lz => xt_rsc_triosy_0_29_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_29_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_28_obj_inst : peaseNTT_core_xt_rsc_triosy_0_28_obj
    PORT MAP(
      xt_rsc_triosy_0_28_lz => xt_rsc_triosy_0_28_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_28_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_27_obj_inst : peaseNTT_core_xt_rsc_triosy_0_27_obj
    PORT MAP(
      xt_rsc_triosy_0_27_lz => xt_rsc_triosy_0_27_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_27_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_26_obj_inst : peaseNTT_core_xt_rsc_triosy_0_26_obj
    PORT MAP(
      xt_rsc_triosy_0_26_lz => xt_rsc_triosy_0_26_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_26_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_25_obj_inst : peaseNTT_core_xt_rsc_triosy_0_25_obj
    PORT MAP(
      xt_rsc_triosy_0_25_lz => xt_rsc_triosy_0_25_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_25_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_24_obj_inst : peaseNTT_core_xt_rsc_triosy_0_24_obj
    PORT MAP(
      xt_rsc_triosy_0_24_lz => xt_rsc_triosy_0_24_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_24_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_23_obj_inst : peaseNTT_core_xt_rsc_triosy_0_23_obj
    PORT MAP(
      xt_rsc_triosy_0_23_lz => xt_rsc_triosy_0_23_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_23_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_22_obj_inst : peaseNTT_core_xt_rsc_triosy_0_22_obj
    PORT MAP(
      xt_rsc_triosy_0_22_lz => xt_rsc_triosy_0_22_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_22_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_21_obj_inst : peaseNTT_core_xt_rsc_triosy_0_21_obj
    PORT MAP(
      xt_rsc_triosy_0_21_lz => xt_rsc_triosy_0_21_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_21_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_20_obj_inst : peaseNTT_core_xt_rsc_triosy_0_20_obj
    PORT MAP(
      xt_rsc_triosy_0_20_lz => xt_rsc_triosy_0_20_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_20_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_19_obj_inst : peaseNTT_core_xt_rsc_triosy_0_19_obj
    PORT MAP(
      xt_rsc_triosy_0_19_lz => xt_rsc_triosy_0_19_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_19_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_18_obj_inst : peaseNTT_core_xt_rsc_triosy_0_18_obj
    PORT MAP(
      xt_rsc_triosy_0_18_lz => xt_rsc_triosy_0_18_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_18_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_17_obj_inst : peaseNTT_core_xt_rsc_triosy_0_17_obj
    PORT MAP(
      xt_rsc_triosy_0_17_lz => xt_rsc_triosy_0_17_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_17_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_16_obj_inst : peaseNTT_core_xt_rsc_triosy_0_16_obj
    PORT MAP(
      xt_rsc_triosy_0_16_lz => xt_rsc_triosy_0_16_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_16_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_15_obj_inst : peaseNTT_core_xt_rsc_triosy_0_15_obj
    PORT MAP(
      xt_rsc_triosy_0_15_lz => xt_rsc_triosy_0_15_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_15_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_14_obj_inst : peaseNTT_core_xt_rsc_triosy_0_14_obj
    PORT MAP(
      xt_rsc_triosy_0_14_lz => xt_rsc_triosy_0_14_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_14_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_13_obj_inst : peaseNTT_core_xt_rsc_triosy_0_13_obj
    PORT MAP(
      xt_rsc_triosy_0_13_lz => xt_rsc_triosy_0_13_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_13_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_12_obj_inst : peaseNTT_core_xt_rsc_triosy_0_12_obj
    PORT MAP(
      xt_rsc_triosy_0_12_lz => xt_rsc_triosy_0_12_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_12_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_11_obj_inst : peaseNTT_core_xt_rsc_triosy_0_11_obj
    PORT MAP(
      xt_rsc_triosy_0_11_lz => xt_rsc_triosy_0_11_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_11_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_10_obj_inst : peaseNTT_core_xt_rsc_triosy_0_10_obj
    PORT MAP(
      xt_rsc_triosy_0_10_lz => xt_rsc_triosy_0_10_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_10_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_9_obj_inst : peaseNTT_core_xt_rsc_triosy_0_9_obj
    PORT MAP(
      xt_rsc_triosy_0_9_lz => xt_rsc_triosy_0_9_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_9_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_8_obj_inst : peaseNTT_core_xt_rsc_triosy_0_8_obj
    PORT MAP(
      xt_rsc_triosy_0_8_lz => xt_rsc_triosy_0_8_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_8_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_7_obj_inst : peaseNTT_core_xt_rsc_triosy_0_7_obj
    PORT MAP(
      xt_rsc_triosy_0_7_lz => xt_rsc_triosy_0_7_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_7_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_6_obj_inst : peaseNTT_core_xt_rsc_triosy_0_6_obj
    PORT MAP(
      xt_rsc_triosy_0_6_lz => xt_rsc_triosy_0_6_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_6_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_5_obj_inst : peaseNTT_core_xt_rsc_triosy_0_5_obj
    PORT MAP(
      xt_rsc_triosy_0_5_lz => xt_rsc_triosy_0_5_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_5_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_4_obj_inst : peaseNTT_core_xt_rsc_triosy_0_4_obj
    PORT MAP(
      xt_rsc_triosy_0_4_lz => xt_rsc_triosy_0_4_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_4_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_3_obj_inst : peaseNTT_core_xt_rsc_triosy_0_3_obj
    PORT MAP(
      xt_rsc_triosy_0_3_lz => xt_rsc_triosy_0_3_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_3_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_2_obj_inst : peaseNTT_core_xt_rsc_triosy_0_2_obj
    PORT MAP(
      xt_rsc_triosy_0_2_lz => xt_rsc_triosy_0_2_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_2_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_1_obj_inst : peaseNTT_core_xt_rsc_triosy_0_1_obj
    PORT MAP(
      xt_rsc_triosy_0_1_lz => xt_rsc_triosy_0_1_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_1_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_xt_rsc_triosy_0_0_obj_inst : peaseNTT_core_xt_rsc_triosy_0_0_obj
    PORT MAP(
      xt_rsc_triosy_0_0_lz => xt_rsc_triosy_0_0_lz,
      core_wten => core_wten,
      xt_rsc_triosy_0_0_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_p_rsc_triosy_obj_inst : peaseNTT_core_p_rsc_triosy_obj
    PORT MAP(
      p_rsc_triosy_lz => p_rsc_triosy_lz,
      core_wten => core_wten,
      p_rsc_triosy_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_r_rsc_triosy_obj_inst : peaseNTT_core_r_rsc_triosy_obj
    PORT MAP(
      r_rsc_triosy_lz => r_rsc_triosy_lz,
      core_wten => core_wten,
      r_rsc_triosy_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_15_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_15_obj
    PORT MAP(
      twiddle_rsc_triosy_0_15_lz => twiddle_rsc_triosy_0_15_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_15_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_14_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_14_obj
    PORT MAP(
      twiddle_rsc_triosy_0_14_lz => twiddle_rsc_triosy_0_14_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_14_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_13_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_13_obj
    PORT MAP(
      twiddle_rsc_triosy_0_13_lz => twiddle_rsc_triosy_0_13_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_13_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_12_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_12_obj
    PORT MAP(
      twiddle_rsc_triosy_0_12_lz => twiddle_rsc_triosy_0_12_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_12_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_11_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_11_obj
    PORT MAP(
      twiddle_rsc_triosy_0_11_lz => twiddle_rsc_triosy_0_11_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_11_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_10_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_10_obj
    PORT MAP(
      twiddle_rsc_triosy_0_10_lz => twiddle_rsc_triosy_0_10_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_10_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_9_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_9_obj
    PORT MAP(
      twiddle_rsc_triosy_0_9_lz => twiddle_rsc_triosy_0_9_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_9_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_8_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_8_obj
    PORT MAP(
      twiddle_rsc_triosy_0_8_lz => twiddle_rsc_triosy_0_8_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_8_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_7_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_7_obj
    PORT MAP(
      twiddle_rsc_triosy_0_7_lz => twiddle_rsc_triosy_0_7_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_7_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_6_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_6_obj
    PORT MAP(
      twiddle_rsc_triosy_0_6_lz => twiddle_rsc_triosy_0_6_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_6_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_5_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_5_obj
    PORT MAP(
      twiddle_rsc_triosy_0_5_lz => twiddle_rsc_triosy_0_5_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_5_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_4_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_4_obj
    PORT MAP(
      twiddle_rsc_triosy_0_4_lz => twiddle_rsc_triosy_0_4_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_4_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_3_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_3_obj
    PORT MAP(
      twiddle_rsc_triosy_0_3_lz => twiddle_rsc_triosy_0_3_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_3_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_2_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_2_obj
    PORT MAP(
      twiddle_rsc_triosy_0_2_lz => twiddle_rsc_triosy_0_2_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_2_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_1_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_1_obj
    PORT MAP(
      twiddle_rsc_triosy_0_1_lz => twiddle_rsc_triosy_0_1_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_1_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_rsc_triosy_0_0_obj_inst : peaseNTT_core_twiddle_rsc_triosy_0_0_obj
    PORT MAP(
      twiddle_rsc_triosy_0_0_lz => twiddle_rsc_triosy_0_0_lz,
      core_wten => core_wten,
      twiddle_rsc_triosy_0_0_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_15_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_15_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_15_lz => twiddle_h_rsc_triosy_0_15_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_15_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_14_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_14_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_14_lz => twiddle_h_rsc_triosy_0_14_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_14_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_13_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_13_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_13_lz => twiddle_h_rsc_triosy_0_13_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_13_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_12_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_12_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_12_lz => twiddle_h_rsc_triosy_0_12_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_12_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_11_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_11_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_11_lz => twiddle_h_rsc_triosy_0_11_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_11_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_10_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_10_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_10_lz => twiddle_h_rsc_triosy_0_10_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_10_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_9_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_9_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_9_lz => twiddle_h_rsc_triosy_0_9_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_9_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_8_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_8_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_8_lz => twiddle_h_rsc_triosy_0_8_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_8_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_7_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_7_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_7_lz => twiddle_h_rsc_triosy_0_7_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_7_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_6_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_6_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_6_lz => twiddle_h_rsc_triosy_0_6_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_6_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_5_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_5_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_5_lz => twiddle_h_rsc_triosy_0_5_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_5_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_4_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_4_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_4_lz => twiddle_h_rsc_triosy_0_4_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_4_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_3_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_3_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_3_lz => twiddle_h_rsc_triosy_0_3_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_3_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_2_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_2_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_2_lz => twiddle_h_rsc_triosy_0_2_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_2_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_1_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_1_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_1_lz => twiddle_h_rsc_triosy_0_1_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_1_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_twiddle_h_rsc_triosy_0_0_obj_inst : peaseNTT_core_twiddle_h_rsc_triosy_0_0_obj
    PORT MAP(
      twiddle_h_rsc_triosy_0_0_lz => twiddle_h_rsc_triosy_0_0_lz,
      core_wten => core_wten,
      twiddle_h_rsc_triosy_0_0_obj_iswt0 => reg_xt_rsc_triosy_1_31_obj_iswt0_cse
    );
  peaseNTT_core_staller_inst : peaseNTT_core_staller
    PORT MAP(
      clk => clk,
      rst => rst,
      core_wen => core_wen,
      core_wten => core_wten,
      twiddle_rsc_0_0_i_wen_comp => twiddle_rsc_0_0_i_wen_comp,
      twiddle_rsc_0_1_i_wen_comp => twiddle_rsc_0_1_i_wen_comp,
      twiddle_rsc_0_2_i_wen_comp => twiddle_rsc_0_2_i_wen_comp,
      twiddle_rsc_0_3_i_wen_comp => twiddle_rsc_0_3_i_wen_comp,
      twiddle_rsc_0_4_i_wen_comp => twiddle_rsc_0_4_i_wen_comp,
      twiddle_rsc_0_5_i_wen_comp => twiddle_rsc_0_5_i_wen_comp,
      twiddle_rsc_0_6_i_wen_comp => twiddle_rsc_0_6_i_wen_comp,
      twiddle_rsc_0_7_i_wen_comp => twiddle_rsc_0_7_i_wen_comp,
      twiddle_rsc_0_8_i_wen_comp => twiddle_rsc_0_8_i_wen_comp,
      twiddle_rsc_0_9_i_wen_comp => twiddle_rsc_0_9_i_wen_comp,
      twiddle_rsc_0_10_i_wen_comp => twiddle_rsc_0_10_i_wen_comp,
      twiddle_rsc_0_11_i_wen_comp => twiddle_rsc_0_11_i_wen_comp,
      twiddle_rsc_0_12_i_wen_comp => twiddle_rsc_0_12_i_wen_comp,
      twiddle_rsc_0_13_i_wen_comp => twiddle_rsc_0_13_i_wen_comp,
      twiddle_rsc_0_14_i_wen_comp => twiddle_rsc_0_14_i_wen_comp,
      twiddle_rsc_0_15_i_wen_comp => twiddle_rsc_0_15_i_wen_comp,
      twiddle_h_rsc_0_0_i_wen_comp => twiddle_h_rsc_0_0_i_wen_comp,
      twiddle_h_rsc_0_1_i_wen_comp => twiddle_h_rsc_0_1_i_wen_comp,
      twiddle_h_rsc_0_2_i_wen_comp => twiddle_h_rsc_0_2_i_wen_comp,
      twiddle_h_rsc_0_3_i_wen_comp => twiddle_h_rsc_0_3_i_wen_comp,
      twiddle_h_rsc_0_4_i_wen_comp => twiddle_h_rsc_0_4_i_wen_comp,
      twiddle_h_rsc_0_5_i_wen_comp => twiddle_h_rsc_0_5_i_wen_comp,
      twiddle_h_rsc_0_6_i_wen_comp => twiddle_h_rsc_0_6_i_wen_comp,
      twiddle_h_rsc_0_7_i_wen_comp => twiddle_h_rsc_0_7_i_wen_comp,
      twiddle_h_rsc_0_8_i_wen_comp => twiddle_h_rsc_0_8_i_wen_comp,
      twiddle_h_rsc_0_9_i_wen_comp => twiddle_h_rsc_0_9_i_wen_comp,
      twiddle_h_rsc_0_10_i_wen_comp => twiddle_h_rsc_0_10_i_wen_comp,
      twiddle_h_rsc_0_11_i_wen_comp => twiddle_h_rsc_0_11_i_wen_comp,
      twiddle_h_rsc_0_12_i_wen_comp => twiddle_h_rsc_0_12_i_wen_comp,
      twiddle_h_rsc_0_13_i_wen_comp => twiddle_h_rsc_0_13_i_wen_comp,
      twiddle_h_rsc_0_14_i_wen_comp => twiddle_h_rsc_0_14_i_wen_comp,
      twiddle_h_rsc_0_15_i_wen_comp => twiddle_h_rsc_0_15_i_wen_comp
    );
  peaseNTT_core_core_fsm_inst : peaseNTT_core_core_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      core_wen => core_wen,
      fsm_output => peaseNTT_core_core_fsm_inst_fsm_output,
      INNER_LOOP1_C_0_tr0 => INNER_LOOP1_nor_tmp,
      INNER_LOOP2_C_0_tr0 => peaseNTT_core_core_fsm_inst_INNER_LOOP2_C_0_tr0,
      INNER_LOOP2_C_0_tr1 => peaseNTT_core_core_fsm_inst_INNER_LOOP2_C_0_tr1,
      INNER_LOOP3_C_0_tr0 => peaseNTT_core_core_fsm_inst_INNER_LOOP3_C_0_tr0,
      INNER_LOOP4_C_0_tr0 => and_dcpl_144,
      INNER_LOOP4_C_0_tr1 => peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1
    );
  fsm_output <= peaseNTT_core_core_fsm_inst_fsm_output;
  peaseNTT_core_core_fsm_inst_INNER_LOOP2_C_0_tr0 <= INNER_LOOP2_nor_tmp AND ((operator_20_false_acc_cse_sva(0))
      XOR (operator_20_false_acc_cse_sva(1)));
  peaseNTT_core_core_fsm_inst_INNER_LOOP2_C_0_tr1 <= NOT INNER_LOOP2_nor_tmp;
  peaseNTT_core_core_fsm_inst_INNER_LOOP3_C_0_tr0 <= NOT(INNER_LOOP3_stage_0 OR INNER_LOOP3_stage_0_2
      OR INNER_LOOP3_stage_0_3 OR INNER_LOOP3_stage_0_4 OR INNER_LOOP3_stage_0_5
      OR INNER_LOOP3_stage_0_6 OR INNER_LOOP3_stage_0_7 OR INNER_LOOP3_stage_0_8
      OR INNER_LOOP3_stage_0_9 OR INNER_LOOP3_stage_0_10 OR INNER_LOOP3_stage_0_11
      OR INNER_LOOP3_stage_0_12);
  peaseNTT_core_core_fsm_inst_INNER_LOOP4_C_0_tr1 <= NOT INNER_LOOP4_nor_tmp;

  or_67_rmff <= ((and_dcpl_147 OR ((NOT INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_191_itm_12)
      AND INNER_LOOP3_stage_0_13)) AND (fsm_output(6))) OR ((and_dcpl_149 OR (INNER_LOOP1_stage_0_13
      AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_160_itm_12))) AND (fsm_output(2)))
      OR and_252_cse OR and_253_cse;
  or_166_rmff <= ((and_dcpl_155 OR (INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_191_itm_12
      AND INNER_LOOP3_stage_0_13)) AND (fsm_output(6))) OR ((and_dcpl_157 OR (INNER_LOOP1_stage_0_13
      AND INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_160_itm_12)) AND (fsm_output(2)))
      OR and_252_cse OR and_253_cse;
  or_248_rmff <= ((and_dcpl_158 OR and_dcpl_147) AND (fsm_output(6))) OR ((and_dcpl_149
      OR and_dcpl_159) AND (fsm_output(2))) OR and_655_cse OR and_656_cse;
  or_347_rmff <= ((and_dcpl_164 OR and_dcpl_155) AND (fsm_output(6))) OR ((and_dcpl_157
      OR and_dcpl_165) AND (fsm_output(2))) OR and_655_cse OR and_656_cse;
  or_429_rmff <= and_1056_cse OR and_1057_cse OR and_1058_cse OR and_1059_cse;
  or_435_rmff <= and_1058_cse OR and_1059_cse;
  or_436_rmff <= and_1056_cse OR and_1057_cse;
  or_512_rmff <= and_1056_cse OR and_1057_cse OR and_1229_cse OR and_1230_cse;
  or_517_rmff <= and_1229_cse OR and_1230_cse;
  or_578_rmff <= and_1363_cse OR and_1364_cse OR and_1058_cse OR and_1059_cse;
  or_584_rmff <= and_1363_cse OR and_1364_cse;
  or_660_rmff <= and_1363_cse OR and_1364_cse OR and_1229_cse OR and_1230_cse;
  and_1665_cse <= INNER_LOOP1_stage_0 AND (fsm_output(2));
  and_1666_cse <= INNER_LOOP2_stage_0 AND (fsm_output(4));
  or_833_rmff <= ((INNER_LOOP3_stage_0_2 OR INNER_LOOP3_stage_0_4 OR INNER_LOOP3_stage_0_3)
      AND (fsm_output(6))) OR ((INNER_LOOP1_stage_0_3 OR INNER_LOOP1_stage_0_2 OR
      INNER_LOOP1_stage_0_4) AND (fsm_output(2))) OR ((INNER_LOOP2_stage_0_3 OR INNER_LOOP2_stage_0_4
      OR INNER_LOOP2_stage_0_2) AND (fsm_output(4))) OR ((INNER_LOOP4_stage_0_2 OR
      INNER_LOOP4_stage_0_4 OR INNER_LOOP4_stage_0_3) AND (fsm_output(8)));
  INNER_LOOP1_tw_h_and_49_cse <= CONV_SL_1_1(operator_33_true_3_lshift_psp_1_0_sva=STD_LOGIC_VECTOR'("00"))
      AND (fsm_output(8));
  INNER_LOOP1_tw_h_and_51_cse <= CONV_SL_1_1(operator_33_true_3_lshift_psp_1_0_sva=STD_LOGIC_VECTOR'("01"))
      AND (fsm_output(8));
  INNER_LOOP1_tw_h_and_53_cse <= CONV_SL_1_1(operator_33_true_3_lshift_psp_1_0_sva=STD_LOGIC_VECTOR'("10"))
      AND (fsm_output(8));
  INNER_LOOP1_tw_h_and_55_cse <= CONV_SL_1_1(operator_33_true_3_lshift_psp_1_0_sva=STD_LOGIC_VECTOR'("11"))
      AND (fsm_output(8));
  INNER_LOOP1_tw_h_and_44_cse <= butterFly2_15_tw_equal_tmp_1 AND (fsm_output(6));
  butterFly2_7_tw_nor_cse <= NOT(CONV_SL_1_1(operator_33_true_2_lshift_psp_2_0_sva(2
      DOWNTO 1)/=STD_LOGIC_VECTOR'("00")));
  INNER_LOOP1_tw_h_and_45_cse <= (operator_33_true_2_lshift_psp_2_0_sva(0)) AND butterFly2_7_tw_nor_cse
      AND (fsm_output(6));
  butterFly2_7_tw_nor_1_cse <= NOT((operator_33_true_2_lshift_psp_2_0_sva(2)) OR
      (operator_33_true_2_lshift_psp_2_0_sva(0)));
  INNER_LOOP1_tw_h_and_46_cse <= (operator_33_true_2_lshift_psp_2_0_sva(1)) AND butterFly2_7_tw_nor_1_cse
      AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_47_cse <= butterFly2_15_tw_equal_tmp_3_1 AND (fsm_output(6));
  butterFly2_7_tw_nor_2_cse <= NOT(CONV_SL_1_1(operator_33_true_2_lshift_psp_2_0_sva(1
      DOWNTO 0)/=STD_LOGIC_VECTOR'("00")));
  INNER_LOOP1_tw_h_and_48_cse <= (operator_33_true_2_lshift_psp_2_0_sva(2)) AND butterFly2_7_tw_nor_2_cse
      AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_50_cse <= butterFly2_15_tw_equal_tmp_5_1 AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_52_cse <= butterFly2_15_tw_equal_tmp_6_1 AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_54_cse <= butterFly2_15_tw_equal_tmp_7_1 AND (fsm_output(6));
  INNER_LOOP1_tw_h_or_9_cse <= INNER_LOOP1_tw_h_and_48_cse OR INNER_LOOP1_tw_h_and_49_cse;
  INNER_LOOP1_tw_h_or_10_cse <= INNER_LOOP1_tw_h_and_50_cse OR INNER_LOOP1_tw_h_and_51_cse;
  INNER_LOOP1_tw_h_or_11_cse <= INNER_LOOP1_tw_h_and_52_cse OR INNER_LOOP1_tw_h_and_53_cse;
  INNER_LOOP1_tw_h_or_12_cse <= INNER_LOOP1_tw_h_and_54_cse OR INNER_LOOP1_tw_h_and_55_cse;
  INNER_LOOP1_tw_h_and_41_cse <= CONV_SL_1_1(operator_33_true_2_lshift_psp_2_0_sva(2
      DOWNTO 1)=STD_LOGIC_VECTOR'("01")) AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_42_cse <= CONV_SL_1_1(operator_33_true_2_lshift_psp_2_0_sva(2
      DOWNTO 1)=STD_LOGIC_VECTOR'("10")) AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_43_cse <= CONV_SL_1_1(operator_33_true_2_lshift_psp_2_0_sva(2
      DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_40_cse <= butterFly2_7_tw_nor_cse AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_37_cse <= (operator_33_true_2_lshift_psp_2_0_sva(0)) AND (NOT
      (operator_33_true_2_lshift_psp_2_0_sva(2))) AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_38_cse <= (operator_33_true_2_lshift_psp_2_0_sva(2)) AND (NOT
      (operator_33_true_2_lshift_psp_2_0_sva(0))) AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_39_cse <= (operator_33_true_2_lshift_psp_2_0_sva(2)) AND (operator_33_true_2_lshift_psp_2_0_sva(0))
      AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_36_cse <= butterFly2_7_tw_nor_1_cse AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_30_cse <= CONV_SL_1_1(operator_33_true_2_lshift_psp_2_0_sva(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("01")) AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_31_cse <= CONV_SL_1_1(operator_33_true_2_lshift_psp_2_0_sva(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("10")) AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_32_cse <= CONV_SL_1_1(operator_33_true_2_lshift_psp_2_0_sva(1
      DOWNTO 0)=STD_LOGIC_VECTOR'("11")) AND (fsm_output(6));
  INNER_LOOP1_tw_h_and_29_cse <= butterFly2_7_tw_nor_2_cse AND (fsm_output(6));
  INNER_LOOP1_tw_h_or_3_cse <= or_dcpl_29 OR INNER_LOOP1_tw_h_and_44_cse;
  INNER_LOOP1_tw_h_or_1_cse <= or_dcpl_29 OR INNER_LOOP1_tw_h_and_36_cse;
  mult_4_t_and_nl <= (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1) AND (fsm_output(2));
  mult_4_t_and_1_nl <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1 AND (fsm_output(2));
  mult_4_t_and_2_nl <= (NOT twiddle_h_rsc_0_0_i_s_raddr_core_4) AND (fsm_output(6));
  mult_4_t_and_3_nl <= twiddle_h_rsc_0_0_i_s_raddr_core_4 AND (fsm_output(6));
  mult_4_t_mux1h_rmff <= MUX1HOT_v_32_6_2(xt_rsc_0_9_i_qa_d_mxwt, xt_rsc_1_9_i_qa_d_mxwt,
      mult_t_mul_cmp_12_a_mx0w3, xt_rsc_0_7_i_qa_d_mxwt, xt_rsc_1_7_i_qa_d_mxwt,
      tmp_23_lpi_3_dfm_mx0, STD_LOGIC_VECTOR'( mult_4_t_and_nl & mult_4_t_and_1_nl
      & (fsm_output(4)) & mult_4_t_and_2_nl & mult_4_t_and_3_nl & (fsm_output(8))));
  INNER_LOOP1_tw_h_or_cse <= or_dcpl_29 OR INNER_LOOP1_tw_h_and_29_cse;
  or_956_rmff <= ((INNER_LOOP3_stage_0_5 OR INNER_LOOP3_stage_0_6 OR INNER_LOOP3_stage_0_7)
      AND (fsm_output(6))) OR ((INNER_LOOP1_stage_0_6 OR INNER_LOOP1_stage_0_7 OR
      INNER_LOOP1_stage_0_5) AND (fsm_output(2))) OR ((INNER_LOOP2_stage_0_6 OR INNER_LOOP2_stage_0_7
      OR INNER_LOOP2_stage_0_5) AND (fsm_output(4))) OR ((INNER_LOOP4_stage_0_5 OR
      INNER_LOOP4_stage_0_6 OR INNER_LOOP4_stage_0_7) AND (fsm_output(8)));
  modulo_add_qelse_and_cse <= core_wen AND INNER_LOOP1_stage_0_11;
  butterFly1_and_cse <= core_wen AND INNER_LOOP1_stage_0_10;
  mult_15_if_and_cse <= core_wen AND INNER_LOOP1_stage_0_9;
  INNER_LOOP1_r_and_7_cse <= core_wen AND INNER_LOOP1_stage_0;
  mult_15_z_and_cse <= core_wen AND INNER_LOOP1_stage_0_8;
  mult_15_z_and_cse_1 <= core_wen AND (INNER_LOOP3_stage_0_8 OR INNER_LOOP2_stage_0_8
      OR INNER_LOOP4_stage_0_8 OR INNER_LOOP1_stage_0_8);
  mult_15_z_and_1_cse <= core_wen AND INNER_LOOP1_stage_0_7;
  mult_15_z_and_2_cse <= core_wen AND INNER_LOOP1_stage_0_6;
  mult_15_z_and_3_cse <= core_wen AND (INNER_LOOP2_stage_0_5 OR INNER_LOOP4_stage_0_5
      OR INNER_LOOP1_stage_0_5 OR INNER_LOOP3_stage_0_5);
  INNER_LOOP1_r_and_20_cse <= core_wen AND INNER_LOOP1_stage_0_5;
  INNER_LOOP1_r_and_23_cse <= core_wen AND INNER_LOOP1_stage_0_4;
  INNER_LOOP1_r_and_26_cse <= core_wen AND INNER_LOOP1_stage_0_3;
  INNER_LOOP1_r_and_29_cse <= core_wen AND INNER_LOOP1_stage_0_2;
  modulo_add_16_qelse_and_cse <= core_wen AND INNER_LOOP2_stage_0_11;
  butterFly1_31_and_cse <= core_wen AND INNER_LOOP2_stage_0_10;
  mult_31_if_and_cse <= core_wen AND INNER_LOOP2_stage_0_9;
  INNER_LOOP2_r_and_3_cse <= core_wen AND INNER_LOOP2_stage_0;
  INNER_LOOP1_r_INNER_LOOP1_r_and_2_cse <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (z_out_33(4 DOWNTO 0)), (fsm_output(4)));
  INNER_LOOP2_r_and_4_cse <= core_wen AND ((fsm_output(3)) OR (INNER_LOOP2_stage_0
      AND (NOT (z_out_33(5))) AND (fsm_output(4))));
  mult_31_z_and_cse <= core_wen AND INNER_LOOP2_stage_0_8;
  mult_31_z_and_1_cse <= core_wen AND INNER_LOOP2_stage_0_7;
  mult_31_z_and_2_cse <= core_wen AND INNER_LOOP2_stage_0_6;
  butterFly1_31_f1_and_4_cse <= core_wen AND INNER_LOOP2_stage_0_5;
  butterFly1_31_f1_and_5_cse <= core_wen AND INNER_LOOP2_stage_0_4;
  butterFly1_31_f1_and_6_cse <= core_wen AND INNER_LOOP2_stage_0_3;
  butterFly1_31_f1_and_7_cse <= core_wen AND (INNER_LOOP4_stage_0_2 OR INNER_LOOP2_stage_0_2);
  c_or_cse <= (fsm_output(4)) OR (fsm_output(8));
  modulo_add_32_qelse_and_cse <= core_wen AND INNER_LOOP3_stage_0_11;
  butterFly2_and_cse <= core_wen AND INNER_LOOP3_stage_0_10;
  mult_47_if_and_cse <= core_wen AND INNER_LOOP3_stage_0_9;
  butterFly2_15_tw_and_cse <= core_wen AND INNER_LOOP3_stage_0;
  INNER_LOOP3_INNER_LOOP3_and_1_cse <= INNER_LOOP3_stage_0 AND (fsm_output(6));
  mult_47_z_and_cse <= core_wen AND INNER_LOOP3_stage_0_8;
  mult_47_z_and_1_cse <= core_wen AND INNER_LOOP3_stage_0_7;
  mult_47_z_and_2_cse <= core_wen AND INNER_LOOP3_stage_0_6;
  INNER_LOOP3_r_and_19_cse <= core_wen AND INNER_LOOP3_stage_0_5;
  INNER_LOOP3_r_and_22_cse <= core_wen AND INNER_LOOP3_stage_0_4;
  INNER_LOOP3_r_and_25_cse <= core_wen AND INNER_LOOP3_stage_0_3;
  INNER_LOOP3_r_and_28_cse <= core_wen AND INNER_LOOP3_stage_0_2;
  modulo_add_48_qelse_and_cse <= core_wen AND INNER_LOOP4_stage_0_11;
  butterFly2_31_and_cse <= core_wen AND INNER_LOOP4_stage_0_10;
  mult_63_if_and_cse <= core_wen AND INNER_LOOP4_stage_0_9;
  INNER_LOOP4_r_and_3_cse <= core_wen AND INNER_LOOP4_stage_0;
  INNER_LOOP1_r_INNER_LOOP1_r_and_6_cse <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"),
      (INNER_LOOP4_r_9_4_sva_2(4 DOWNTO 0)), (fsm_output(8)));
  INNER_LOOP4_INNER_LOOP4_and_1_cse <= INNER_LOOP4_stage_0 AND (fsm_output(8));
  INNER_LOOP4_r_and_4_cse <= core_wen AND ((fsm_output(7)) OR (INNER_LOOP4_stage_0
      AND (NOT (INNER_LOOP4_r_9_4_sva_2(5))) AND (fsm_output(8))));
  mult_63_z_and_cse <= core_wen AND INNER_LOOP4_stage_0_8;
  mult_63_z_and_1_cse <= core_wen AND INNER_LOOP4_stage_0_7;
  mult_63_z_and_2_cse <= core_wen AND INNER_LOOP4_stage_0_6;
  butterFly2_31_f1_and_4_cse <= core_wen AND INNER_LOOP4_stage_0_5;
  butterFly2_31_f1_and_5_cse <= core_wen AND INNER_LOOP4_stage_0_4;
  butterFly2_31_f1_and_6_cse <= core_wen AND INNER_LOOP4_stage_0_3;
  mult_t_mul_cmp_a_mx0w2 <= MUX_v_32_2_2(xt_rsc_0_31_i_qa_d_mxwt, xt_rsc_1_31_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_1_a_mx0w0 <= MUX_v_32_2_2(xt_rsc_0_31_i_qa_d_mxwt, xt_rsc_1_31_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  mult_t_mul_cmp_2_a_mx0w2 <= MUX_v_32_2_2(xt_rsc_0_27_i_qa_d_mxwt, xt_rsc_1_27_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_4_a_mx0w2 <= MUX_v_32_2_2(xt_rsc_0_23_i_qa_d_mxwt, xt_rsc_1_23_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_5_a_mx0w2 <= MUX_v_32_2_2(xt_rsc_0_21_i_qa_d_mxwt, xt_rsc_1_21_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_12_a_mx0w3 <= MUX_v_32_2_2(yt_rsc_0_9_i_qa_d, yt_rsc_1_9_i_qa_d,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_6_a_mx0w2 <= MUX_v_32_2_2(xt_rsc_0_19_i_qa_d_mxwt, xt_rsc_1_19_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_11_a_mx0w3 <= MUX_v_32_2_2(yt_rsc_0_11_i_qa_d, yt_rsc_1_11_i_qa_d,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_7_a_mx0w2 <= MUX_v_32_2_2(xt_rsc_0_17_i_qa_d_mxwt, xt_rsc_1_17_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_10_a_mx0w3 <= MUX_v_32_2_2(yt_rsc_0_13_i_qa_d, yt_rsc_1_13_i_qa_d,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_8_a_mx0w2 <= MUX_v_32_2_2(xt_rsc_0_15_i_qa_d_mxwt, xt_rsc_1_15_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_9_a_mx0w3 <= MUX_v_32_2_2(yt_rsc_0_15_i_qa_d, yt_rsc_1_15_i_qa_d,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_9_a_mx0w0 <= MUX_v_32_2_2(xt_rsc_0_15_i_qa_d_mxwt, xt_rsc_1_15_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  mult_t_mul_cmp_9_a_mx0w2 <= MUX_v_32_2_2(xt_rsc_0_13_i_qa_d_mxwt, xt_rsc_1_13_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_10_a_mx0w0 <= MUX_v_32_2_2(xt_rsc_0_13_i_qa_d_mxwt, xt_rsc_1_13_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  mult_t_mul_cmp_10_a_mx0w2 <= MUX_v_32_2_2(xt_rsc_0_11_i_qa_d_mxwt, xt_rsc_1_11_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_11_a_mx0w0 <= MUX_v_32_2_2(xt_rsc_0_11_i_qa_d_mxwt, xt_rsc_1_11_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  mult_t_mul_cmp_11_a_mx0w2 <= MUX_v_32_2_2(xt_rsc_0_9_i_qa_d_mxwt, xt_rsc_1_9_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_13_a_mx0w0 <= MUX_v_32_2_2(xt_rsc_0_7_i_qa_d_mxwt, xt_rsc_1_7_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  mult_t_mul_cmp_13_a_mx0w2 <= MUX_v_32_2_2(xt_rsc_0_5_i_qa_d_mxwt, xt_rsc_1_5_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_14_a_mx0w0 <= MUX_v_32_2_2(xt_rsc_0_5_i_qa_d_mxwt, xt_rsc_1_5_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  mult_t_mul_cmp_14_a_mx0w2 <= MUX_v_32_2_2(xt_rsc_0_3_i_qa_d_mxwt, xt_rsc_1_3_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_t_mul_cmp_15_a_mx0w0 <= MUX_v_32_2_2(xt_rsc_0_3_i_qa_d_mxwt, xt_rsc_1_3_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  mult_t_mul_cmp_15_a_mx0w2 <= MUX_v_32_2_2(xt_rsc_0_1_i_qa_d_mxwt, xt_rsc_1_1_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  operator_20_false_acc_cse_sva_mx0w0 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(butterFly2_19_tw_asn_itm
      & c_1_sva) + UNSIGNED'( "111"), 3));
  mult_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_z_asn_itm_4) - UNSIGNED(reg_mult_z_asn_itm_1_cse),
      32));
  mult_1_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_1_z_asn_itm_4)
      - UNSIGNED(reg_mult_1_z_asn_itm_1_cse), 32));
  mult_2_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_2_z_asn_itm_4)
      - UNSIGNED(reg_mult_2_z_asn_itm_1_cse), 32));
  mult_3_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_3_z_asn_itm_4)
      - UNSIGNED(reg_mult_3_z_asn_itm_1_cse), 32));
  mult_4_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_4_z_asn_itm_4)
      - UNSIGNED(reg_mult_4_z_asn_itm_1_cse), 32));
  mult_5_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_5_z_asn_itm_4)
      - UNSIGNED(reg_mult_5_z_asn_itm_1_cse), 32));
  mult_6_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_6_z_asn_itm_4)
      - UNSIGNED(reg_mult_6_z_asn_itm_1_cse), 32));
  mult_7_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_7_z_asn_itm_4)
      - UNSIGNED(reg_mult_7_z_asn_itm_1_cse), 32));
  mult_8_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_8_z_asn_itm_4)
      - UNSIGNED(reg_mult_8_z_asn_itm_1_cse), 32));
  mult_9_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_9_z_asn_itm_4)
      - UNSIGNED(reg_mult_9_z_asn_itm_1_cse), 32));
  mult_10_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_10_z_asn_itm_4)
      - UNSIGNED(reg_mult_10_z_asn_itm_1_cse), 32));
  mult_11_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_11_z_asn_itm_4)
      - UNSIGNED(reg_mult_11_z_asn_itm_1_cse), 32));
  mult_12_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_12_z_asn_itm_4)
      - UNSIGNED(reg_mult_12_z_asn_itm_1_cse), 32));
  mult_13_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_13_z_asn_itm_4)
      - UNSIGNED(reg_mult_13_z_asn_itm_1_cse), 32));
  mult_14_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_14_z_asn_itm_4)
      - UNSIGNED(reg_mult_14_z_asn_itm_1_cse), 32));
  mult_15_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_15_z_asn_itm_4)
      - UNSIGNED(reg_mult_15_z_asn_itm_1_cse), 32));
  tmp_93_lpi_3_dfm_mx0 <= MUX_v_32_2_2(xt_rsc_0_29_i_qa_d_mxwt, xt_rsc_1_29_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  tmp_91_lpi_3_dfm_mx0 <= MUX_v_32_2_2(xt_rsc_0_27_i_qa_d_mxwt, xt_rsc_1_27_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  tmp_89_lpi_3_dfm_mx0 <= MUX_v_32_2_2(xt_rsc_0_25_i_qa_d_mxwt, xt_rsc_1_25_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  tmp_87_lpi_3_dfm_mx0 <= MUX_v_32_2_2(xt_rsc_0_23_i_qa_d_mxwt, xt_rsc_1_23_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  tmp_85_lpi_3_dfm_mx0 <= MUX_v_32_2_2(xt_rsc_0_21_i_qa_d_mxwt, xt_rsc_1_21_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  tmp_83_lpi_3_dfm_mx0 <= MUX_v_32_2_2(xt_rsc_0_19_i_qa_d_mxwt, xt_rsc_1_19_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  tmp_81_lpi_3_dfm_mx0 <= MUX_v_32_2_2(xt_rsc_0_17_i_qa_d_mxwt, xt_rsc_1_17_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  tmp_65_lpi_3_dfm_mx0 <= MUX_v_32_2_2(xt_rsc_0_1_i_qa_d_mxwt, xt_rsc_1_1_i_qa_d_mxwt,
      INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
  INNER_LOOP1_r_9_4_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(INNER_LOOP1_r_9_4_sva_4_0),
      5), 6) + UNSIGNED'( "000001"), 6));
  INNER_LOOP1_tw_and_psp_sva_1 <= operator_33_true_return_8_4_sva AND INNER_LOOP1_r_9_4_sva_4_0;
  mult_15_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_34, mult_15_res_sva_1, mult_15_slc_32_svs_st_1);
  mult_14_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_35, mult_14_res_sva_1, mult_14_slc_32_svs_st_1);
  mult_13_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_36, mult_13_res_sva_1, mult_13_slc_32_svs_st_1);
  mult_12_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_51, mult_12_res_sva_1, mult_12_slc_32_svs_st_1);
  mult_11_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_63, mult_11_res_sva_1, mult_11_slc_32_svs_st_1);
  mult_10_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_38, mult_10_res_sva_1, mult_10_slc_32_svs_st_1);
  mult_9_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_61, mult_9_res_sva_1, mult_9_slc_32_svs_st_1);
  mult_8_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_59, mult_8_res_sva_1, mult_8_slc_32_svs_st_1);
  mult_7_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_57, mult_7_res_sva_1, mult_7_slc_32_svs_st_1);
  mult_6_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_53, mult_6_res_sva_1, mult_6_slc_32_svs_st_1);
  mult_5_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_103, mult_5_res_sva_1, mult_5_slc_32_svs_st_1);
  mult_4_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_108, mult_4_res_sva_1, mult_4_slc_32_svs_st_1);
  mult_3_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_104, mult_3_res_sva_1, mult_3_slc_32_svs_st_1);
  mult_2_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_107, mult_2_res_sva_1, mult_2_slc_32_svs_st_1);
  mult_1_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_109, mult_1_res_sva_1, mult_1_slc_32_svs_st_1);
  mult_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_105, mult_res_sva_1, mult_slc_32_svs_st_1);
  mult_25_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_25_z_asn_itm_4)
      - UNSIGNED(reg_mult_9_z_asn_itm_1_cse), 32));
  mult_26_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_26_z_asn_itm_4)
      - UNSIGNED(reg_mult_10_z_asn_itm_1_cse), 32));
  mult_27_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_27_z_asn_itm_4)
      - UNSIGNED(reg_mult_11_z_asn_itm_1_cse), 32));
  mult_28_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_28_z_asn_itm_4)
      - UNSIGNED(reg_mult_12_z_asn_itm_1_cse), 32));
  mult_29_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_29_z_asn_itm_4)
      - UNSIGNED(reg_mult_13_z_asn_itm_1_cse), 32));
  mult_30_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_30_z_asn_itm_4)
      - UNSIGNED(reg_mult_14_z_asn_itm_1_cse), 32));
  mult_31_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_31_z_asn_itm_4)
      - UNSIGNED(reg_mult_15_z_asn_itm_1_cse), 32));
  tmp_31_lpi_3_dfm_mx0 <= MUX_v_32_2_2(yt_rsc_0_31_i_qa_d, yt_rsc_1_31_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
  tmp_29_lpi_3_dfm_mx0 <= MUX_v_32_2_2(yt_rsc_0_29_i_qa_d, yt_rsc_1_29_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
  tmp_27_lpi_3_dfm_mx0 <= MUX_v_32_2_2(yt_rsc_0_27_i_qa_d, yt_rsc_1_27_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
  tmp_25_lpi_3_dfm_mx0 <= MUX_v_32_2_2(yt_rsc_0_25_i_qa_d, yt_rsc_1_25_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
  tmp_23_lpi_3_dfm_mx0 <= MUX_v_32_2_2(yt_rsc_0_23_i_qa_d, yt_rsc_1_23_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
  tmp_21_lpi_3_dfm_mx0 <= MUX_v_32_2_2(yt_rsc_0_21_i_qa_d, yt_rsc_1_21_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
  tmp_19_lpi_3_dfm_mx0 <= MUX_v_32_2_2(yt_rsc_0_19_i_qa_d, yt_rsc_1_19_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
  tmp_17_lpi_3_dfm_mx0 <= MUX_v_32_2_2(yt_rsc_0_17_i_qa_d, yt_rsc_1_17_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
  tmp_7_lpi_3_dfm_mx0 <= MUX_v_32_2_2(yt_rsc_0_7_i_qa_d, yt_rsc_1_7_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
  tmp_5_lpi_3_dfm_mx0 <= MUX_v_32_2_2(yt_rsc_0_5_i_qa_d, yt_rsc_1_5_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
  tmp_3_lpi_3_dfm_mx0 <= MUX_v_32_2_2(yt_rsc_0_3_i_qa_d, yt_rsc_1_3_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
  tmp_1_lpi_3_dfm_mx0 <= MUX_v_32_2_2(yt_rsc_0_1_i_qa_d, yt_rsc_1_1_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_31_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_51, mult_31_res_sva_1, mult_31_slc_32_svs_st_1);
  mult_30_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_34, mult_30_res_sva_1, mult_30_slc_32_svs_st_1);
  mult_29_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_57, mult_29_res_sva_1, mult_29_slc_32_svs_st_1);
  mult_28_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_63, mult_28_res_sva_1, mult_28_slc_32_svs_st_1);
  mult_27_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_53, mult_27_res_sva_1, mult_27_slc_32_svs_st_1);
  mult_26_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_36, mult_26_res_sva_1, mult_26_slc_32_svs_st_1);
  mult_25_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_35, mult_25_res_sva_1, mult_25_slc_32_svs_st_1);
  mult_24_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_59, mult_24_res_sva_1, mult_24_slc_32_svs_st_1);
  mult_23_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_61, mult_23_res_sva_1, mult_23_slc_32_svs_st_1);
  mult_22_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_22_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_22_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_22_if_acc_nl),
      32)), mult_22_res_sva_1, mult_22_slc_32_svs_st_1);
  mult_21_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_21_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_21_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_21_if_acc_nl),
      32)), mult_21_res_sva_1, mult_21_slc_32_svs_st_1);
  mult_20_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_20_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_20_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_20_if_acc_nl),
      32)), mult_20_res_sva_1, mult_20_slc_32_svs_st_1);
  mult_19_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_19_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_19_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_19_if_acc_nl),
      32)), mult_19_res_sva_1, mult_19_slc_32_svs_st_1);
  mult_18_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_18_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_18_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_18_if_acc_nl),
      32)), mult_18_res_sva_1, mult_18_slc_32_svs_st_1);
  mult_17_if_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_17_res_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_17_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_17_if_acc_nl),
      32)), mult_17_res_sva_1, mult_17_slc_32_svs_st_1);
  mult_16_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_106, mult_16_res_sva_1, mult_16_slc_32_svs_st_1);
  mult_32_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_32_z_asn_itm_4)
      - UNSIGNED(reg_mult_z_asn_itm_1_cse), 32));
  mult_33_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_33_z_asn_itm_4)
      - UNSIGNED(reg_mult_5_z_asn_itm_1_cse), 32));
  mult_34_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_34_z_asn_itm_4)
      - UNSIGNED(reg_mult_8_z_asn_itm_1_cse), 32));
  mult_35_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_35_z_asn_itm_4)
      - UNSIGNED(reg_mult_13_z_asn_itm_1_cse), 32));
  mult_36_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_36_z_asn_itm_4)
      - UNSIGNED(reg_mult_15_z_asn_itm_1_cse), 32));
  mult_37_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_37_z_asn_itm_4)
      - UNSIGNED(reg_mult_11_z_asn_itm_1_cse), 32));
  mult_38_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_38_z_asn_itm_4)
      - UNSIGNED(reg_mult_7_z_asn_itm_1_cse), 32));
  mult_39_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_39_z_asn_itm_4)
      - UNSIGNED(reg_mult_3_z_asn_itm_1_cse), 32));
  mult_40_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_40_z_asn_itm_4)
      - UNSIGNED(reg_mult_2_z_asn_itm_1_cse), 32));
  mult_41_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_41_z_asn_itm_4)
      - UNSIGNED(reg_mult_10_z_asn_itm_1_cse), 32));
  mult_42_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_42_z_asn_itm_4)
      - UNSIGNED(reg_mult_14_z_asn_itm_1_cse), 32));
  mult_43_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_43_z_asn_itm_4)
      - UNSIGNED(reg_mult_6_z_asn_itm_1_cse), 32));
  mult_44_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_44_z_asn_itm_4)
      - UNSIGNED(reg_mult_4_z_asn_itm_1_cse), 32));
  mult_45_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_45_z_asn_itm_4)
      - UNSIGNED(reg_mult_12_z_asn_itm_1_cse), 32));
  mult_46_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_46_z_asn_itm_4)
      - UNSIGNED(reg_mult_9_z_asn_itm_1_cse), 32));
  mult_47_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_47_z_asn_itm_4)
      - UNSIGNED(reg_mult_1_z_asn_itm_1_cse), 32));
  tmp_125_lpi_3_dfm_mx0 <= MUX_v_32_2_2(xt_rsc_0_29_i_qa_d_mxwt, xt_rsc_1_29_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  tmp_121_lpi_3_dfm_mx0 <= MUX_v_32_2_2(xt_rsc_0_25_i_qa_d_mxwt, xt_rsc_1_25_i_qa_d_mxwt,
      twiddle_h_rsc_0_0_i_s_raddr_core_4);
  mult_47_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_51, mult_47_res_sva_1, mult_47_slc_32_svs_st_1);
  mult_46_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_105, mult_46_res_sva_1, mult_46_slc_32_svs_st_1);
  mult_45_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_107, mult_45_res_sva_1, mult_45_slc_32_svs_st_1);
  mult_44_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_106, mult_44_res_sva_1, mult_44_slc_32_svs_st_1);
  mult_43_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_102, mult_43_res_sva_1, mult_43_slc_32_svs_st_1);
  mult_42_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_108, mult_42_res_sva_1, mult_42_slc_32_svs_st_1);
  mult_41_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_103, mult_41_res_sva_1, mult_41_slc_32_svs_st_1);
  mult_40_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_109, mult_40_res_sva_1, mult_40_slc_32_svs_st_1);
  mult_39_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_104, mult_39_res_sva_1, mult_39_slc_32_svs_st_1);
  mult_38_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_96, mult_38_res_sva_1, mult_38_slc_32_svs_st_1);
  mult_37_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_95, mult_37_res_sva_1, mult_37_slc_32_svs_st_1);
  mult_36_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_94, mult_36_res_sva_1, mult_36_slc_32_svs_st_1);
  mult_35_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_93, mult_35_res_sva_1, mult_35_slc_32_svs_st_1);
  mult_34_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_92, mult_34_res_sva_1, mult_34_slc_32_svs_st_1);
  mult_33_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_88, mult_33_res_sva_1, mult_33_slc_32_svs_st_1);
  mult_32_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_87, mult_32_res_sva_1, mult_32_slc_32_svs_st_1);
  mult_48_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_48_z_asn_itm_4)
      - UNSIGNED(reg_mult_1_z_asn_itm_1_cse), 32));
  mult_49_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_49_z_asn_itm_4)
      - UNSIGNED(reg_mult_9_z_asn_itm_1_cse), 32));
  mult_50_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_50_z_asn_itm_4)
      - UNSIGNED(reg_mult_12_z_asn_itm_1_cse), 32));
  mult_51_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_51_z_asn_itm_4)
      - UNSIGNED(reg_mult_4_z_asn_itm_1_cse), 32));
  mult_52_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_52_z_asn_itm_4)
      - UNSIGNED(reg_mult_6_z_asn_itm_1_cse), 32));
  mult_53_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_53_z_asn_itm_4)
      - UNSIGNED(reg_mult_14_z_asn_itm_1_cse), 32));
  mult_54_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_54_z_asn_itm_4)
      - UNSIGNED(reg_mult_10_z_asn_itm_1_cse), 32));
  mult_55_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_55_z_asn_itm_4)
      - UNSIGNED(reg_mult_2_z_asn_itm_1_cse), 32));
  mult_56_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_56_z_asn_itm_4)
      - UNSIGNED(reg_mult_3_z_asn_itm_1_cse), 32));
  mult_57_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_57_z_asn_itm_4)
      - UNSIGNED(reg_mult_7_z_asn_itm_1_cse), 32));
  mult_58_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_58_z_asn_itm_4)
      - UNSIGNED(reg_mult_11_z_asn_itm_1_cse), 32));
  mult_59_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_59_z_asn_itm_4)
      - UNSIGNED(reg_mult_15_z_asn_itm_1_cse), 32));
  mult_60_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_60_z_asn_itm_4)
      - UNSIGNED(reg_mult_13_z_asn_itm_1_cse), 32));
  mult_61_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_61_z_asn_itm_4)
      - UNSIGNED(reg_mult_8_z_asn_itm_1_cse), 32));
  mult_62_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_62_z_asn_itm_4)
      - UNSIGNED(reg_mult_5_z_asn_itm_1_cse), 32));
  mult_63_res_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_63_z_asn_itm_4)
      - UNSIGNED(reg_mult_z_asn_itm_1_cse), 32));
  INNER_LOOP4_r_9_4_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(INNER_LOOP4_r_9_4_sva_4_0),
      5), 6) + UNSIGNED'( "000001"), 6));
  mult_63_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_107, mult_63_res_sva_1, mult_63_slc_32_svs_st_1);
  mult_62_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_105, mult_62_res_sva_1, mult_62_slc_32_svs_st_1);
  mult_61_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_104, mult_61_res_sva_1, mult_61_slc_32_svs_st_1);
  mult_60_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_103, mult_60_res_sva_1, mult_60_slc_32_svs_st_1);
  mult_59_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_102, mult_59_res_sva_1, mult_59_slc_32_svs_st_1);
  mult_58_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_100, mult_58_res_sva_1, mult_58_slc_32_svs_st_1);
  mult_57_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_99, mult_57_res_sva_1, mult_57_slc_32_svs_st_1);
  mult_56_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_98, mult_56_res_sva_1, mult_56_slc_32_svs_st_1);
  mult_55_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_97, mult_55_res_sva_1, mult_55_slc_32_svs_st_1);
  mult_54_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_96, mult_54_res_sva_1, mult_54_slc_32_svs_st_1);
  mult_53_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_95, mult_53_res_sva_1, mult_53_slc_32_svs_st_1);
  mult_52_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_94, mult_52_res_sva_1, mult_52_slc_32_svs_st_1);
  mult_51_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_93, mult_51_res_sva_1, mult_51_slc_32_svs_st_1);
  mult_50_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_92, mult_50_res_sva_1, mult_50_slc_32_svs_st_1);
  mult_49_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_88, mult_49_res_sva_1, mult_49_slc_32_svs_st_1);
  mult_48_res_lpi_3_dfm_mx0 <= MUX_v_32_2_2(z_out_87, mult_48_res_sva_1, mult_48_slc_32_svs_st_1);
  INNER_LOOP4_nor_tmp <= NOT(INNER_LOOP4_stage_0 OR INNER_LOOP4_stage_0_2 OR INNER_LOOP4_stage_0_3
      OR INNER_LOOP4_stage_0_4 OR INNER_LOOP4_stage_0_5 OR INNER_LOOP4_stage_0_6
      OR INNER_LOOP4_stage_0_7 OR INNER_LOOP4_stage_0_8 OR INNER_LOOP4_stage_0_9
      OR INNER_LOOP4_stage_0_10 OR INNER_LOOP4_stage_0_11 OR INNER_LOOP4_stage_0_12);
  INNER_LOOP2_nor_tmp <= NOT(INNER_LOOP2_stage_0 OR INNER_LOOP2_stage_0_2 OR INNER_LOOP2_stage_0_3
      OR INNER_LOOP2_stage_0_4 OR INNER_LOOP2_stage_0_5 OR INNER_LOOP2_stage_0_6
      OR INNER_LOOP2_stage_0_7 OR INNER_LOOP2_stage_0_8 OR INNER_LOOP2_stage_0_9
      OR INNER_LOOP2_stage_0_10 OR INNER_LOOP2_stage_0_11 OR INNER_LOOP2_stage_0_12);
  INNER_LOOP1_nor_tmp <= NOT(INNER_LOOP1_stage_0 OR INNER_LOOP1_stage_0_2 OR INNER_LOOP1_stage_0_3
      OR INNER_LOOP1_stage_0_4 OR INNER_LOOP1_stage_0_5 OR INNER_LOOP1_stage_0_6
      OR INNER_LOOP1_stage_0_7 OR INNER_LOOP1_stage_0_8 OR INNER_LOOP1_stage_0_9
      OR INNER_LOOP1_stage_0_10 OR INNER_LOOP1_stage_0_11 OR INNER_LOOP1_stage_0_12);
  and_dcpl_144 <= INNER_LOOP4_nor_tmp AND c_1_sva_1;
  and_dcpl_147 <= INNER_LOOP3_stage_0_12 AND (NOT INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_11);
  and_dcpl_149 <= INNER_LOOP1_stage_0_12 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_11);
  and_dcpl_151 <= INNER_LOOP2_stage_0 AND (NOT (INNER_LOOP2_r_9_4_sva_4_0(4)));
  and_dcpl_153 <= INNER_LOOP4_stage_0 AND (NOT (INNER_LOOP4_r_9_4_sva_4_0(4)));
  and_dcpl_155 <= INNER_LOOP3_stage_0_12 AND INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_11;
  and_dcpl_157 <= INNER_LOOP1_stage_0_12 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_11;
  and_dcpl_158 <= (NOT INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_10) AND INNER_LOOP3_stage_0_11;
  and_dcpl_159 <= INNER_LOOP1_stage_0_11 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_10);
  and_dcpl_161 <= INNER_LOOP2_stage_0 AND (INNER_LOOP2_r_9_4_sva_4_0(4));
  and_dcpl_163 <= INNER_LOOP4_stage_0 AND (INNER_LOOP4_r_9_4_sva_4_0(4));
  and_dcpl_164 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_10 AND INNER_LOOP3_stage_0_11;
  and_dcpl_165 <= INNER_LOOP1_stage_0_11 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_10;
  and_dcpl_174 <= INNER_LOOP3_stage_0 AND (operator_33_true_2_lshift_psp_2_0_sva(0));
  and_dcpl_175 <= INNER_LOOP4_stage_0 AND (operator_33_true_3_lshift_psp_1_0_sva(0));
  and_dcpl_176 <= INNER_LOOP3_stage_0 AND (operator_33_true_2_lshift_psp_2_0_sva(1));
  or_dcpl_29 <= (fsm_output(2)) OR (fsm_output(4));
  and_252_cse <= (and_dcpl_151 OR ((NOT INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4302_itm_1)
      AND INNER_LOOP2_stage_0_2)) AND (fsm_output(4));
  and_253_cse <= (and_dcpl_153 OR (INNER_LOOP4_stage_0_2 AND (NOT INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4377_itm_1)))
      AND (fsm_output(8));
  and_655_cse <= (and_dcpl_161 OR (INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4302_itm_1
      AND INNER_LOOP2_stage_0_2)) AND (fsm_output(4));
  and_656_cse <= (and_dcpl_163 OR (INNER_LOOP4_stage_0_2 AND INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4377_itm_1))
      AND (fsm_output(8));
  and_1058_cse <= INNER_LOOP2_stage_0_12 AND (NOT INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_11)
      AND (fsm_output(4));
  and_1059_cse <= INNER_LOOP4_stage_0_12 AND (NOT INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_11)
      AND (fsm_output(8));
  and_1056_cse <= INNER_LOOP3_stage_0 AND (NOT (INNER_LOOP3_r_9_4_sva_4_0(4))) AND
      (fsm_output(6));
  and_1057_cse <= INNER_LOOP1_stage_0 AND (NOT (INNER_LOOP1_r_9_4_sva_4_0(4))) AND
      (fsm_output(2));
  and_1229_cse <= INNER_LOOP2_stage_0_12 AND INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_11
      AND (fsm_output(4));
  and_1230_cse <= INNER_LOOP4_stage_0_12 AND INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_11
      AND (fsm_output(8));
  and_1363_cse <= INNER_LOOP3_stage_0 AND (INNER_LOOP3_r_9_4_sva_4_0(4)) AND (fsm_output(6));
  and_1364_cse <= INNER_LOOP1_stage_0 AND (INNER_LOOP1_r_9_4_sva_4_0(4)) AND (fsm_output(2));
  and_1686_cse <= and_dcpl_175 AND (fsm_output(8));
  and_1695_cse <= INNER_LOOP4_stage_0 AND (operator_33_true_3_lshift_psp_1_0_sva(1))
      AND (fsm_output(8));
  and_1704_cse <= and_dcpl_175 AND (operator_33_true_3_lshift_psp_1_0_sva(1)) AND
      (fsm_output(8));
  and_1929_cse <= (NOT (operator_33_true_3_lshift_psp_1_0_sva(0))) AND (fsm_output(8));
  or_tmp_804 <= or_dcpl_29 OR and_1929_cse;
  or_tmp_806 <= (operator_33_true_3_lshift_psp_1_0_sva(0)) AND (fsm_output(8));
  and_1944_cse <= (NOT (operator_33_true_3_lshift_psp_1_0_sva(1))) AND (fsm_output(8));
  or_tmp_812 <= (operator_33_true_2_lshift_psp_2_0_sva(2)) AND (fsm_output(6));
  and_1948_cse <= (NOT (operator_33_true_2_lshift_psp_2_0_sva(2))) AND (fsm_output(6));
  or_tmp_814 <= (operator_33_true_3_lshift_psp_1_0_sva(1)) AND (fsm_output(8));
  or_tmp_827 <= (operator_33_true_2_lshift_psp_2_0_sva(1)) AND (fsm_output(6));
  and_1978_cse <= (NOT (operator_33_true_2_lshift_psp_2_0_sva(1))) AND (fsm_output(6));
  or_tmp_835 <= (operator_33_true_2_lshift_psp_2_0_sva(0)) AND (fsm_output(6));
  and_1994_cse <= (NOT (operator_33_true_2_lshift_psp_2_0_sva(0))) AND (fsm_output(6));
  or_tmp_888 <= and_1978_cse OR or_dcpl_29;
  or_tmp_895 <= and_1994_cse OR or_dcpl_29;
  butterFly1_and_ssc <= NOT((modulo_sub_base_sva_1(31)) OR (fsm_output(6)));
  butterFly1_and_ssc_2 <= (NOT (modulo_sub_base_32_sva_1(31))) AND (fsm_output(6));
  butterFly1_and_ssc_3 <= (modulo_sub_base_32_sva_1(31)) AND (fsm_output(6));
  butterFly1_1_and_ssc <= NOT((modulo_sub_base_1_sva_1(31)) OR (fsm_output(6)));
  butterFly1_1_and_ssc_2 <= (NOT (modulo_sub_base_33_sva_1(31))) AND (fsm_output(6));
  butterFly1_1_and_ssc_3 <= (modulo_sub_base_33_sva_1(31)) AND (fsm_output(6));
  butterFly1_2_and_ssc <= NOT((modulo_sub_base_2_sva_1(31)) OR (fsm_output(6)));
  butterFly1_2_and_ssc_2 <= (NOT (modulo_sub_base_34_sva_1(31))) AND (fsm_output(6));
  butterFly1_2_and_ssc_3 <= (modulo_sub_base_34_sva_1(31)) AND (fsm_output(6));
  butterFly1_3_and_ssc <= NOT((modulo_sub_base_3_sva_1(31)) OR (fsm_output(6)));
  butterFly1_3_and_ssc_2 <= (NOT (modulo_sub_base_35_sva_1(31))) AND (fsm_output(6));
  butterFly1_3_and_ssc_3 <= (modulo_sub_base_35_sva_1(31)) AND (fsm_output(6));
  butterFly1_4_and_ssc <= NOT((modulo_sub_base_4_sva_1(31)) OR (fsm_output(6)));
  butterFly1_4_and_ssc_2 <= (NOT (modulo_sub_base_36_sva_1(31))) AND (fsm_output(6));
  butterFly1_4_and_ssc_3 <= (modulo_sub_base_36_sva_1(31)) AND (fsm_output(6));
  butterFly1_5_and_ssc <= NOT((modulo_sub_base_5_sva_1(31)) OR (fsm_output(6)));
  butterFly1_5_and_ssc_2 <= (NOT (modulo_sub_base_37_sva_1(31))) AND (fsm_output(6));
  butterFly1_5_and_ssc_3 <= (modulo_sub_base_37_sva_1(31)) AND (fsm_output(6));
  butterFly1_6_and_ssc <= NOT((modulo_sub_base_6_sva_1(31)) OR (fsm_output(6)));
  butterFly1_6_and_ssc_2 <= (NOT (modulo_sub_base_38_sva_1(31))) AND (fsm_output(6));
  butterFly1_6_and_ssc_3 <= (modulo_sub_base_38_sva_1(31)) AND (fsm_output(6));
  butterFly1_7_and_ssc <= NOT((modulo_sub_base_7_sva_1(31)) OR (fsm_output(6)));
  butterFly1_7_and_ssc_2 <= (NOT (modulo_sub_base_39_sva_1(31))) AND (fsm_output(6));
  butterFly1_7_and_ssc_3 <= (modulo_sub_base_39_sva_1(31)) AND (fsm_output(6));
  butterFly1_8_and_ssc <= NOT((modulo_sub_base_8_sva_1(31)) OR (fsm_output(6)));
  butterFly1_8_and_ssc_2 <= (NOT (modulo_sub_base_40_sva_1(31))) AND (fsm_output(6));
  butterFly1_8_and_ssc_3 <= (modulo_sub_base_40_sva_1(31)) AND (fsm_output(6));
  butterFly1_9_and_ssc <= NOT((modulo_sub_base_9_sva_1(31)) OR (fsm_output(6)));
  butterFly1_9_and_ssc_2 <= (NOT (modulo_sub_base_41_sva_1(31))) AND (fsm_output(6));
  butterFly1_9_and_ssc_3 <= (modulo_sub_base_41_sva_1(31)) AND (fsm_output(6));
  butterFly1_10_and_ssc <= NOT((modulo_sub_base_10_sva_1(31)) OR (fsm_output(6)));
  butterFly1_10_and_ssc_2 <= (NOT (modulo_sub_base_42_sva_1(31))) AND (fsm_output(6));
  butterFly1_10_and_ssc_3 <= (modulo_sub_base_42_sva_1(31)) AND (fsm_output(6));
  butterFly1_11_and_ssc <= NOT((modulo_sub_base_11_sva_1(31)) OR (fsm_output(6)));
  butterFly1_11_and_ssc_2 <= (NOT (modulo_sub_base_43_sva_1(31))) AND (fsm_output(6));
  butterFly1_11_and_ssc_3 <= (modulo_sub_base_43_sva_1(31)) AND (fsm_output(6));
  butterFly1_12_and_ssc <= NOT((modulo_sub_base_12_sva_1(31)) OR (fsm_output(6)));
  butterFly1_12_and_ssc_2 <= (NOT (modulo_sub_base_44_sva_1(31))) AND (fsm_output(6));
  butterFly1_12_and_ssc_3 <= (modulo_sub_base_44_sva_1(31)) AND (fsm_output(6));
  butterFly1_13_and_ssc <= NOT((modulo_sub_base_13_sva_1(31)) OR (fsm_output(6)));
  butterFly1_13_and_ssc_2 <= (NOT (modulo_sub_base_45_sva_1(31))) AND (fsm_output(6));
  butterFly1_13_and_ssc_3 <= (modulo_sub_base_45_sva_1(31)) AND (fsm_output(6));
  butterFly1_14_and_ssc <= NOT((modulo_sub_base_14_sva_1(31)) OR (fsm_output(6)));
  butterFly1_14_and_ssc_2 <= (NOT (modulo_sub_base_46_sva_1(31))) AND (fsm_output(6));
  butterFly1_14_and_ssc_3 <= (modulo_sub_base_46_sva_1(31)) AND (fsm_output(6));
  butterFly1_15_and_ssc <= NOT((modulo_sub_base_15_sva_1(31)) OR (fsm_output(6)));
  butterFly1_15_and_ssc_2 <= (NOT (modulo_sub_base_47_sva_1(31))) AND (fsm_output(6));
  butterFly1_15_and_ssc_3 <= (modulo_sub_base_47_sva_1(31)) AND (fsm_output(6));
  butterFly1_mux_nl <= MUX_s_1_2_2((z_out_81(31)), (z_out_80(31)), butterFly1_and_ssc_3);
  butterFly1_and_4_rmff <= butterFly1_mux_nl AND (NOT(butterFly1_and_ssc OR butterFly1_and_ssc_2));
  butterFly1_and_1_nl <= (modulo_sub_base_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_sva_1(30 DOWNTO 0)),
      (z_out_81(30 DOWNTO 0)), (modulo_sub_base_32_sva_1(30 DOWNTO 0)), (z_out_80(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_and_ssc & butterFly1_and_1_nl & butterFly1_and_ssc_2
      & butterFly1_and_ssc_3));
  butterFly1_1_mux_nl <= MUX_s_1_2_2((z_out_79(31)), (z_out_78(31)), butterFly1_1_and_ssc_3);
  butterFly1_1_and_4_rmff <= butterFly1_1_mux_nl AND (NOT(butterFly1_1_and_ssc OR
      butterFly1_1_and_ssc_2));
  butterFly1_1_and_1_nl <= (modulo_sub_base_1_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_1_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_1_sva_1(30 DOWNTO
      0)), (z_out_79(30 DOWNTO 0)), (modulo_sub_base_33_sva_1(30 DOWNTO 0)), (z_out_78(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_1_and_ssc & butterFly1_1_and_1_nl
      & butterFly1_1_and_ssc_2 & butterFly1_1_and_ssc_3));
  butterFly1_2_mux_nl <= MUX_s_1_2_2((z_out_77(31)), (z_out_76(31)), butterFly1_2_and_ssc_3);
  butterFly1_2_and_4_rmff <= butterFly1_2_mux_nl AND (NOT(butterFly1_2_and_ssc OR
      butterFly1_2_and_ssc_2));
  butterFly1_2_and_1_nl <= (modulo_sub_base_2_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_2_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_2_sva_1(30 DOWNTO
      0)), (z_out_77(30 DOWNTO 0)), (modulo_sub_base_34_sva_1(30 DOWNTO 0)), (z_out_76(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_2_and_ssc & butterFly1_2_and_1_nl
      & butterFly1_2_and_ssc_2 & butterFly1_2_and_ssc_3));
  butterFly1_3_mux_nl <= MUX_s_1_2_2((z_out_75(31)), (z_out_74(31)), butterFly1_3_and_ssc_3);
  butterFly1_3_and_4_rmff <= butterFly1_3_mux_nl AND (NOT(butterFly1_3_and_ssc OR
      butterFly1_3_and_ssc_2));
  butterFly1_3_and_1_nl <= (modulo_sub_base_3_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_3_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_3_sva_1(30 DOWNTO
      0)), (z_out_75(30 DOWNTO 0)), (modulo_sub_base_35_sva_1(30 DOWNTO 0)), (z_out_74(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_3_and_ssc & butterFly1_3_and_1_nl
      & butterFly1_3_and_ssc_2 & butterFly1_3_and_ssc_3));
  butterFly1_4_mux_nl <= MUX_s_1_2_2((z_out_73(31)), (z_out_72(31)), butterFly1_4_and_ssc_3);
  butterFly1_4_and_4_rmff <= butterFly1_4_mux_nl AND (NOT(butterFly1_4_and_ssc OR
      butterFly1_4_and_ssc_2));
  butterFly1_4_and_1_nl <= (modulo_sub_base_4_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_4_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_4_sva_1(30 DOWNTO
      0)), (z_out_73(30 DOWNTO 0)), (modulo_sub_base_36_sva_1(30 DOWNTO 0)), (z_out_72(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_4_and_ssc & butterFly1_4_and_1_nl
      & butterFly1_4_and_ssc_2 & butterFly1_4_and_ssc_3));
  butterFly1_5_mux_nl <= MUX_s_1_2_2((z_out_71(31)), (z_out_70(31)), butterFly1_5_and_ssc_3);
  butterFly1_5_and_4_rmff <= butterFly1_5_mux_nl AND (NOT(butterFly1_5_and_ssc OR
      butterFly1_5_and_ssc_2));
  butterFly1_5_and_1_nl <= (modulo_sub_base_5_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_5_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_5_sva_1(30 DOWNTO
      0)), (z_out_71(30 DOWNTO 0)), (modulo_sub_base_37_sva_1(30 DOWNTO 0)), (z_out_70(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_5_and_ssc & butterFly1_5_and_1_nl
      & butterFly1_5_and_ssc_2 & butterFly1_5_and_ssc_3));
  butterFly1_6_mux_nl <= MUX_s_1_2_2((z_out_69(31)), (z_out_68(31)), butterFly1_6_and_ssc_3);
  butterFly1_6_and_4_rmff <= butterFly1_6_mux_nl AND (NOT(butterFly1_6_and_ssc OR
      butterFly1_6_and_ssc_2));
  butterFly1_6_and_1_nl <= (modulo_sub_base_6_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_6_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_6_sva_1(30 DOWNTO
      0)), (z_out_69(30 DOWNTO 0)), (modulo_sub_base_38_sva_1(30 DOWNTO 0)), (z_out_68(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_6_and_ssc & butterFly1_6_and_1_nl
      & butterFly1_6_and_ssc_2 & butterFly1_6_and_ssc_3));
  butterFly1_7_mux_nl <= MUX_s_1_2_2((z_out_67(31)), (z_out_66(31)), butterFly1_7_and_ssc_3);
  butterFly1_7_and_4_rmff <= butterFly1_7_mux_nl AND (NOT(butterFly1_7_and_ssc OR
      butterFly1_7_and_ssc_2));
  butterFly1_7_and_1_nl <= (modulo_sub_base_7_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_7_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_7_sva_1(30 DOWNTO
      0)), (z_out_67(30 DOWNTO 0)), (modulo_sub_base_39_sva_1(30 DOWNTO 0)), (z_out_66(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_7_and_ssc & butterFly1_7_and_1_nl
      & butterFly1_7_and_ssc_2 & butterFly1_7_and_ssc_3));
  butterFly1_8_mux_nl <= MUX_s_1_2_2((z_out_65(31)), (z_out_64(31)), butterFly1_8_and_ssc_3);
  butterFly1_8_and_4_rmff <= butterFly1_8_mux_nl AND (NOT(butterFly1_8_and_ssc OR
      butterFly1_8_and_ssc_2));
  butterFly1_8_and_1_nl <= (modulo_sub_base_8_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_8_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_8_sva_1(30 DOWNTO
      0)), (z_out_65(30 DOWNTO 0)), (modulo_sub_base_40_sva_1(30 DOWNTO 0)), (z_out_64(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_8_and_ssc & butterFly1_8_and_1_nl
      & butterFly1_8_and_ssc_2 & butterFly1_8_and_ssc_3));
  butterFly1_9_mux_nl <= MUX_s_1_2_2((z_out_49(31)), (z_out_62(31)), butterFly1_9_and_ssc_3);
  butterFly1_9_and_4_rmff <= butterFly1_9_mux_nl AND (NOT(butterFly1_9_and_ssc OR
      butterFly1_9_and_ssc_2));
  butterFly1_9_and_1_nl <= (modulo_sub_base_9_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_9_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_9_sva_1(30 DOWNTO
      0)), (z_out_49(30 DOWNTO 0)), (modulo_sub_base_41_sva_1(30 DOWNTO 0)), (z_out_62(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_9_and_ssc & butterFly1_9_and_1_nl
      & butterFly1_9_and_ssc_2 & butterFly1_9_and_ssc_3));
  butterFly1_10_mux_nl <= MUX_s_1_2_2((z_out_47(31)), (z_out_60(31)), butterFly1_10_and_ssc_3);
  butterFly1_10_and_4_rmff <= butterFly1_10_mux_nl AND (NOT(butterFly1_10_and_ssc
      OR butterFly1_10_and_ssc_2));
  butterFly1_10_and_1_nl <= (modulo_sub_base_10_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_10_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_10_sva_1(30 DOWNTO
      0)), (z_out_47(30 DOWNTO 0)), (modulo_sub_base_42_sva_1(30 DOWNTO 0)), (z_out_60(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_10_and_ssc & butterFly1_10_and_1_nl
      & butterFly1_10_and_ssc_2 & butterFly1_10_and_ssc_3));
  butterFly1_11_mux_nl <= MUX_s_1_2_2((z_out_45(31)), (z_out_58(31)), butterFly1_11_and_ssc_3);
  butterFly1_11_and_4_rmff <= butterFly1_11_mux_nl AND (NOT(butterFly1_11_and_ssc
      OR butterFly1_11_and_ssc_2));
  butterFly1_11_and_1_nl <= (modulo_sub_base_11_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_11_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_11_sva_1(30 DOWNTO
      0)), (z_out_45(30 DOWNTO 0)), (modulo_sub_base_43_sva_1(30 DOWNTO 0)), (z_out_58(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_11_and_ssc & butterFly1_11_and_1_nl
      & butterFly1_11_and_ssc_2 & butterFly1_11_and_ssc_3));
  butterFly1_12_mux_nl <= MUX_s_1_2_2((z_out_43(31)), (z_out_56(31)), butterFly1_12_and_ssc_3);
  butterFly1_12_and_4_rmff <= butterFly1_12_mux_nl AND (NOT(butterFly1_12_and_ssc
      OR butterFly1_12_and_ssc_2));
  butterFly1_12_and_1_nl <= (modulo_sub_base_12_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_12_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_12_sva_1(30 DOWNTO
      0)), (z_out_43(30 DOWNTO 0)), (modulo_sub_base_44_sva_1(30 DOWNTO 0)), (z_out_56(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_12_and_ssc & butterFly1_12_and_1_nl
      & butterFly1_12_and_ssc_2 & butterFly1_12_and_ssc_3));
  butterFly1_13_mux_nl <= MUX_s_1_2_2((z_out_41(31)), (z_out_54(31)), butterFly1_13_and_ssc_3);
  butterFly1_13_and_4_rmff <= butterFly1_13_mux_nl AND (NOT(butterFly1_13_and_ssc
      OR butterFly1_13_and_ssc_2));
  butterFly1_13_and_1_nl <= (modulo_sub_base_13_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_13_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_13_sva_1(30 DOWNTO
      0)), (z_out_41(30 DOWNTO 0)), (modulo_sub_base_45_sva_1(30 DOWNTO 0)), (z_out_54(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_13_and_ssc & butterFly1_13_and_1_nl
      & butterFly1_13_and_ssc_2 & butterFly1_13_and_ssc_3));
  butterFly1_14_mux_nl <= MUX_s_1_2_2((z_out_39(31)), (z_out_52(31)), butterFly1_14_and_ssc_3);
  butterFly1_14_and_4_rmff <= butterFly1_14_mux_nl AND (NOT(butterFly1_14_and_ssc
      OR butterFly1_14_and_ssc_2));
  butterFly1_14_and_1_nl <= (modulo_sub_base_14_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_14_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_14_sva_1(30 DOWNTO
      0)), (z_out_39(30 DOWNTO 0)), (modulo_sub_base_46_sva_1(30 DOWNTO 0)), (z_out_52(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_14_and_ssc & butterFly1_14_and_1_nl
      & butterFly1_14_and_ssc_2 & butterFly1_14_and_ssc_3));
  butterFly1_15_mux_nl <= MUX_s_1_2_2((z_out_37(31)), (z_out_50(31)), butterFly1_15_and_ssc_3);
  butterFly1_15_and_4_rmff <= butterFly1_15_mux_nl AND (NOT(butterFly1_15_and_ssc
      OR butterFly1_15_and_ssc_2));
  butterFly1_15_and_1_nl <= (modulo_sub_base_15_sva_1(31)) AND (NOT (fsm_output(6)));
  butterFly1_15_mux1h_2_rmff <= MUX1HOT_v_31_4_2((modulo_sub_base_15_sva_1(30 DOWNTO
      0)), (z_out_37(30 DOWNTO 0)), (modulo_sub_base_47_sva_1(30 DOWNTO 0)), (z_out_50(30
      DOWNTO 0)), STD_LOGIC_VECTOR'( butterFly1_15_and_ssc & butterFly1_15_and_1_nl
      & butterFly1_15_and_ssc_2 & butterFly1_15_and_ssc_3));
  yt_rsc_0_0_i_adra_d_pff <= MUX1HOT_v_4_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_290_itm_11,
      (INNER_LOOP2_r_9_4_sva_4_0(3 DOWNTO 0)), INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_321_itm_11,
      (INNER_LOOP4_r_9_4_sva_4_0(3 DOWNTO 0)), STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  yt_rsc_0_0_i_da_d_pff <= MUX_v_32_2_2(modulo_add_qr_lpi_3_dfm_1, modulo_add_32_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_0_i_wea_d_pff <= (and_dcpl_147 AND (fsm_output(6))) OR (and_dcpl_149 AND
      (fsm_output(2)));
  yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff <= (and_dcpl_151 AND (fsm_output(4)))
      OR (and_dcpl_153 AND (fsm_output(8)));
  yt_rsc_0_1_i_da_d_pff <= MUX_v_32_2_2(modulo_add_1_qr_lpi_3_dfm_1, modulo_add_33_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_2_i_da_d_pff <= MUX_v_32_2_2(modulo_add_2_qr_lpi_3_dfm_1, modulo_add_34_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_3_i_da_d_pff <= MUX_v_32_2_2(modulo_add_3_qr_lpi_3_dfm_1, modulo_add_35_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_4_i_da_d_pff <= MUX_v_32_2_2(modulo_add_4_qr_lpi_3_dfm_1, modulo_add_36_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_5_i_da_d_pff <= MUX_v_32_2_2(modulo_add_5_qr_lpi_3_dfm_1, modulo_add_37_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_6_i_da_d_pff <= MUX_v_32_2_2(modulo_add_6_qr_lpi_3_dfm_1, modulo_add_38_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_7_i_da_d_pff <= MUX_v_32_2_2(modulo_add_7_qr_lpi_3_dfm_1, modulo_add_39_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_8_i_da_d_pff <= MUX_v_32_2_2(modulo_add_8_qr_lpi_3_dfm_1, modulo_add_40_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_9_i_da_d_pff <= MUX_v_32_2_2(modulo_add_9_qr_lpi_3_dfm_1, modulo_add_41_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_10_i_da_d_pff <= MUX_v_32_2_2(modulo_add_10_qr_lpi_3_dfm_1, modulo_add_42_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_11_i_da_d_pff <= MUX_v_32_2_2(modulo_add_11_qr_lpi_3_dfm_1, modulo_add_43_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_12_i_da_d_pff <= MUX_v_32_2_2(modulo_add_12_qr_lpi_3_dfm_1, modulo_add_44_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_13_i_da_d_pff <= MUX_v_32_2_2(modulo_add_13_qr_lpi_3_dfm_1, modulo_add_45_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_14_i_da_d_pff <= MUX_v_32_2_2(modulo_add_14_qr_lpi_3_dfm_1, modulo_add_46_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_15_i_da_d_pff <= MUX_v_32_2_2(modulo_add_15_qr_lpi_3_dfm_1, modulo_add_47_qr_lpi_3_dfm_1,
      fsm_output(6));
  yt_rsc_0_16_i_adra_d_pff <= MUX1HOT_v_4_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_306_itm_11,
      (INNER_LOOP2_r_9_4_sva_4_0(3 DOWNTO 0)), INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_337_itm_11,
      (INNER_LOOP4_r_9_4_sva_4_0(3 DOWNTO 0)), STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  yt_rsc_0_16_i_wea_d_pff <= (and_dcpl_155 AND (fsm_output(6))) OR (and_dcpl_157
      AND (fsm_output(2)));
  yt_rsc_1_0_i_adra_d_pff <= MUX1HOT_v_4_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_385_itm_10,
      (INNER_LOOP2_r_9_4_sva_4_0(3 DOWNTO 0)), INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_416_itm_10,
      (INNER_LOOP4_r_9_4_sva_4_0(3 DOWNTO 0)), STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  yt_rsc_1_0_i_da_d <= butterFly1_and_4_rmff & butterFly1_mux1h_2_rmff;
  yt_rsc_1_0_i_wea_d_pff <= (and_dcpl_158 AND (fsm_output(6))) OR (and_dcpl_159 AND
      (fsm_output(2)));
  yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff <= (and_dcpl_161 AND (fsm_output(4)))
      OR (and_dcpl_163 AND (fsm_output(8)));
  yt_rsc_1_1_i_da_d <= butterFly1_1_and_4_rmff & butterFly1_1_mux1h_2_rmff;
  yt_rsc_1_2_i_da_d <= butterFly1_2_and_4_rmff & butterFly1_2_mux1h_2_rmff;
  yt_rsc_1_3_i_da_d <= butterFly1_3_and_4_rmff & butterFly1_3_mux1h_2_rmff;
  yt_rsc_1_4_i_da_d <= butterFly1_4_and_4_rmff & butterFly1_4_mux1h_2_rmff;
  yt_rsc_1_5_i_da_d <= butterFly1_5_and_4_rmff & butterFly1_5_mux1h_2_rmff;
  yt_rsc_1_6_i_da_d <= butterFly1_6_and_4_rmff & butterFly1_6_mux1h_2_rmff;
  yt_rsc_1_7_i_da_d <= butterFly1_7_and_4_rmff & butterFly1_7_mux1h_2_rmff;
  yt_rsc_1_8_i_da_d <= butterFly1_8_and_4_rmff & butterFly1_8_mux1h_2_rmff;
  yt_rsc_1_9_i_da_d <= butterFly1_9_and_4_rmff & butterFly1_9_mux1h_2_rmff;
  yt_rsc_1_10_i_da_d <= butterFly1_10_and_4_rmff & butterFly1_10_mux1h_2_rmff;
  yt_rsc_1_11_i_da_d <= butterFly1_11_and_4_rmff & butterFly1_11_mux1h_2_rmff;
  yt_rsc_1_12_i_da_d <= butterFly1_12_and_4_rmff & butterFly1_12_mux1h_2_rmff;
  yt_rsc_1_13_i_da_d <= butterFly1_13_and_4_rmff & butterFly1_13_mux1h_2_rmff;
  yt_rsc_1_14_i_da_d <= butterFly1_14_and_4_rmff & butterFly1_14_mux1h_2_rmff;
  yt_rsc_1_15_i_da_d <= butterFly1_15_and_4_rmff & butterFly1_15_mux1h_2_rmff;
  yt_rsc_1_16_i_adra_d_pff <= MUX1HOT_v_4_4_2(INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_401_itm_10,
      (INNER_LOOP2_r_9_4_sva_4_0(3 DOWNTO 0)), INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_432_itm_10,
      (INNER_LOOP4_r_9_4_sva_4_0(3 DOWNTO 0)), STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  yt_rsc_1_16_i_da_d <= butterFly1_and_4_rmff & butterFly1_mux1h_2_rmff;
  yt_rsc_1_16_i_wea_d_pff <= (and_dcpl_164 AND (fsm_output(6))) OR (and_dcpl_165
      AND (fsm_output(2)));
  yt_rsc_1_17_i_da_d <= butterFly1_1_and_4_rmff & butterFly1_1_mux1h_2_rmff;
  yt_rsc_1_18_i_da_d <= butterFly1_2_and_4_rmff & butterFly1_2_mux1h_2_rmff;
  yt_rsc_1_19_i_da_d <= butterFly1_3_and_4_rmff & butterFly1_3_mux1h_2_rmff;
  yt_rsc_1_20_i_da_d <= butterFly1_4_and_4_rmff & butterFly1_4_mux1h_2_rmff;
  yt_rsc_1_21_i_da_d <= butterFly1_5_and_4_rmff & butterFly1_5_mux1h_2_rmff;
  yt_rsc_1_22_i_da_d <= butterFly1_6_and_4_rmff & butterFly1_6_mux1h_2_rmff;
  yt_rsc_1_23_i_da_d <= butterFly1_7_and_4_rmff & butterFly1_7_mux1h_2_rmff;
  yt_rsc_1_24_i_da_d <= butterFly1_8_and_4_rmff & butterFly1_8_mux1h_2_rmff;
  yt_rsc_1_25_i_da_d <= butterFly1_9_and_4_rmff & butterFly1_9_mux1h_2_rmff;
  yt_rsc_1_26_i_da_d <= butterFly1_10_and_4_rmff & butterFly1_10_mux1h_2_rmff;
  yt_rsc_1_27_i_da_d <= butterFly1_11_and_4_rmff & butterFly1_11_mux1h_2_rmff;
  yt_rsc_1_28_i_da_d <= butterFly1_12_and_4_rmff & butterFly1_12_mux1h_2_rmff;
  yt_rsc_1_29_i_da_d <= butterFly1_13_and_4_rmff & butterFly1_13_mux1h_2_rmff;
  yt_rsc_1_30_i_da_d <= butterFly1_14_and_4_rmff & butterFly1_14_mux1h_2_rmff;
  yt_rsc_1_31_i_da_d <= butterFly1_15_and_4_rmff & butterFly1_15_mux1h_2_rmff;
  xt_rsc_0_0_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_9_4_sva_4_0(3 DOWNTO
      0)), INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_290_itm_11, (INNER_LOOP3_r_9_4_sva_4_0(3
      DOWNTO 0)), INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_321_itm_11, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  xt_rsc_0_0_i_da_d_pff <= MUX_v_32_2_2(modulo_add_16_qr_lpi_3_dfm_1, modulo_add_48_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_0_i_wea_d_pff <= xt_rsc_0_0_i_wea_d_iff;
  xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_1_i_da_d_pff <= MUX_v_32_2_2(modulo_add_17_qr_lpi_3_dfm_1, modulo_add_49_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_1_i_wea_d_pff <= xt_rsc_0_1_i_wea_d_iff;
  xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_2_i_da_d_pff <= MUX_v_32_2_2(modulo_add_18_qr_lpi_3_dfm_1, modulo_add_50_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_2_i_wea_d_pff <= xt_rsc_0_2_i_wea_d_iff;
  xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_3_i_da_d_pff <= MUX_v_32_2_2(modulo_add_19_qr_lpi_3_dfm_1, modulo_add_51_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_3_i_wea_d_pff <= xt_rsc_0_3_i_wea_d_iff;
  xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_4_i_da_d_pff <= MUX_v_32_2_2(modulo_add_20_qr_lpi_3_dfm_1, modulo_add_52_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_4_i_wea_d_pff <= xt_rsc_0_4_i_wea_d_iff;
  xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_5_i_da_d_pff <= MUX_v_32_2_2(modulo_add_21_qr_lpi_3_dfm_1, modulo_add_53_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_5_i_wea_d_pff <= xt_rsc_0_5_i_wea_d_iff;
  xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_6_i_da_d_pff <= MUX_v_32_2_2(modulo_add_22_qr_lpi_3_dfm_1, modulo_add_54_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_6_i_wea_d_pff <= xt_rsc_0_6_i_wea_d_iff;
  xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_7_i_da_d_pff <= MUX_v_32_2_2(modulo_add_23_qr_lpi_3_dfm_1, modulo_add_55_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_7_i_wea_d_pff <= xt_rsc_0_7_i_wea_d_iff;
  xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_8_i_da_d_pff <= MUX_v_32_2_2(modulo_add_24_qr_lpi_3_dfm_1, modulo_add_56_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_8_i_wea_d_pff <= xt_rsc_0_8_i_wea_d_iff;
  xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_9_i_da_d_pff <= MUX_v_32_2_2(modulo_add_25_qr_lpi_3_dfm_1, modulo_add_57_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_9_i_wea_d_pff <= xt_rsc_0_9_i_wea_d_iff;
  xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_10_i_da_d_pff <= MUX_v_32_2_2(modulo_add_26_qr_lpi_3_dfm_1, modulo_add_58_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_10_i_wea_d_pff <= xt_rsc_0_10_i_wea_d_iff;
  xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_11_i_da_d_pff <= MUX_v_32_2_2(modulo_add_27_qr_lpi_3_dfm_1, modulo_add_59_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_11_i_wea_d_pff <= xt_rsc_0_11_i_wea_d_iff;
  xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_12_i_da_d_pff <= MUX_v_32_2_2(modulo_add_28_qr_lpi_3_dfm_1, modulo_add_60_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_12_i_wea_d_pff <= xt_rsc_0_12_i_wea_d_iff;
  xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_13_i_da_d_pff <= MUX_v_32_2_2(modulo_add_29_qr_lpi_3_dfm_1, modulo_add_61_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_13_i_wea_d_pff <= xt_rsc_0_13_i_wea_d_iff;
  xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_14_i_da_d_pff <= MUX_v_32_2_2(modulo_add_30_qr_lpi_3_dfm_1, modulo_add_62_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_14_i_wea_d_pff <= xt_rsc_0_14_i_wea_d_iff;
  xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_15_i_da_d_pff <= MUX_v_32_2_2(modulo_add_31_qr_lpi_3_dfm_1, modulo_add_63_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_0_15_i_wea_d_pff <= xt_rsc_0_15_i_wea_d_iff;
  xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_16_i_adra_d_pff <= MUX1HOT_v_4_4_2((INNER_LOOP1_r_9_4_sva_4_0(3 DOWNTO
      0)), INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_306_itm_11, (INNER_LOOP3_r_9_4_sva_4_0(3
      DOWNTO 0)), INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_337_itm_11, STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  xt_rsc_0_16_i_wea_d_pff <= xt_rsc_0_16_i_wea_d_iff;
  xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_17_i_wea_d_pff <= xt_rsc_0_17_i_wea_d_iff;
  xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_18_i_wea_d_pff <= xt_rsc_0_18_i_wea_d_iff;
  xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_19_i_wea_d_pff <= xt_rsc_0_19_i_wea_d_iff;
  xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_20_i_wea_d_pff <= xt_rsc_0_20_i_wea_d_iff;
  xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_21_i_wea_d_pff <= xt_rsc_0_21_i_wea_d_iff;
  xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_22_i_wea_d_pff <= xt_rsc_0_22_i_wea_d_iff;
  xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_23_i_wea_d_pff <= xt_rsc_0_23_i_wea_d_iff;
  xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_24_i_wea_d_pff <= xt_rsc_0_24_i_wea_d_iff;
  xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_25_i_wea_d_pff <= xt_rsc_0_25_i_wea_d_iff;
  xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_26_i_wea_d_pff <= xt_rsc_0_26_i_wea_d_iff;
  xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_27_i_wea_d_pff <= xt_rsc_0_27_i_wea_d_iff;
  xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_28_i_wea_d_pff <= xt_rsc_0_28_i_wea_d_iff;
  xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_29_i_wea_d_pff <= xt_rsc_0_29_i_wea_d_iff;
  xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_30_i_wea_d_pff <= xt_rsc_0_30_i_wea_d_iff;
  xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_0_31_i_wea_d_pff <= xt_rsc_0_31_i_wea_d_iff;
  xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_0_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_16_qr_lpi_3_dfm_1, modulo_sub_48_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_0_i_wea_d_pff <= xt_rsc_1_0_i_wea_d_iff;
  xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_1_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_17_qr_lpi_3_dfm_1, modulo_sub_49_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_1_i_wea_d_pff <= xt_rsc_1_1_i_wea_d_iff;
  xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_2_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_18_qr_lpi_3_dfm_1, modulo_sub_50_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_2_i_wea_d_pff <= xt_rsc_1_2_i_wea_d_iff;
  xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_3_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_19_qr_lpi_3_dfm_1, modulo_sub_51_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_3_i_wea_d_pff <= xt_rsc_1_3_i_wea_d_iff;
  xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_4_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_20_qr_lpi_3_dfm_1, modulo_sub_52_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_4_i_wea_d_pff <= xt_rsc_1_4_i_wea_d_iff;
  xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_5_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_21_qr_lpi_3_dfm_1, modulo_sub_53_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_5_i_wea_d_pff <= xt_rsc_1_5_i_wea_d_iff;
  xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_6_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_22_qr_lpi_3_dfm_1, modulo_sub_54_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_6_i_wea_d_pff <= xt_rsc_1_6_i_wea_d_iff;
  xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_7_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_23_qr_lpi_3_dfm_1, modulo_sub_55_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_7_i_wea_d_pff <= xt_rsc_1_7_i_wea_d_iff;
  xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_8_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_24_qr_lpi_3_dfm_1, modulo_sub_56_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_8_i_wea_d_pff <= xt_rsc_1_8_i_wea_d_iff;
  xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_9_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_25_qr_lpi_3_dfm_1, modulo_sub_57_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_9_i_wea_d_pff <= xt_rsc_1_9_i_wea_d_iff;
  xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_10_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_26_qr_lpi_3_dfm_1, modulo_sub_58_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_10_i_wea_d_pff <= xt_rsc_1_10_i_wea_d_iff;
  xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_11_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_27_qr_lpi_3_dfm_1, modulo_sub_59_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_11_i_wea_d_pff <= xt_rsc_1_11_i_wea_d_iff;
  xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_12_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_28_qr_lpi_3_dfm_1, modulo_sub_60_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_12_i_wea_d_pff <= xt_rsc_1_12_i_wea_d_iff;
  xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_13_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_29_qr_lpi_3_dfm_1, modulo_sub_61_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_13_i_wea_d_pff <= xt_rsc_1_13_i_wea_d_iff;
  xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_14_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_30_qr_lpi_3_dfm_1, modulo_sub_62_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_14_i_wea_d_pff <= xt_rsc_1_14_i_wea_d_iff;
  xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_15_i_da_d_pff <= MUX_v_32_2_2(modulo_sub_31_qr_lpi_3_dfm_1, modulo_sub_63_qr_lpi_3_dfm_1,
      fsm_output(8));
  xt_rsc_1_15_i_wea_d_pff <= xt_rsc_1_15_i_wea_d_iff;
  xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_16_i_wea_d_pff <= xt_rsc_1_16_i_wea_d_iff;
  xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_17_i_wea_d_pff <= xt_rsc_1_17_i_wea_d_iff;
  xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_18_i_wea_d_pff <= xt_rsc_1_18_i_wea_d_iff;
  xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_19_i_wea_d_pff <= xt_rsc_1_19_i_wea_d_iff;
  xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_20_i_wea_d_pff <= xt_rsc_1_20_i_wea_d_iff;
  xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_21_i_wea_d_pff <= xt_rsc_1_21_i_wea_d_iff;
  xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_22_i_wea_d_pff <= xt_rsc_1_22_i_wea_d_iff;
  xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_23_i_wea_d_pff <= xt_rsc_1_23_i_wea_d_iff;
  xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_24_i_wea_d_pff <= xt_rsc_1_24_i_wea_d_iff;
  xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_25_i_wea_d_pff <= xt_rsc_1_25_i_wea_d_iff;
  xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_26_i_wea_d_pff <= xt_rsc_1_26_i_wea_d_iff;
  xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_27_i_wea_d_pff <= xt_rsc_1_27_i_wea_d_iff;
  xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_28_i_wea_d_pff <= xt_rsc_1_28_i_wea_d_iff;
  xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_29_i_wea_d_pff <= xt_rsc_1_29_i_wea_d_iff;
  xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_30_i_wea_d_pff <= xt_rsc_1_30_i_wea_d_iff;
  xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  xt_rsc_1_31_i_wea_d_pff <= xt_rsc_1_31_i_wea_d_iff;
  xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d <= xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d_reg;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND ((fsm_output(9)) OR (fsm_output(0)))) = '1' ) THEN
        p_sva <= p_rsci_idat;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( core_wen = '1' ) THEN
        c_1_sva <= (operator_20_false_acc_cse_sva(0)) OR (NOT (fsm_output(4)));
        reg_twiddle_rsc_0_0_i_s_raddr_core_3_0_cse <= MUX1HOT_v_4_4_2((INNER_LOOP1_tw_and_psp_sva_1(3
            DOWNTO 0)), INNER_LOOP2_tw_and_nl, (INNER_LOOP3_r_9_4_sva_4_0(3 DOWNTO
            0)), (INNER_LOOP4_r_9_4_sva_4_0(3 DOWNTO 0)), STD_LOGIC_VECTOR'( (fsm_output(2))
            & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
        reg_twiddle_rsc_0_1_i_s_raddr_core_4_0_cse <= MUX_v_5_2_2(INNER_LOOP3_r_9_4_sva_4_0,
            INNER_LOOP4_r_9_4_sva_4_0, fsm_output(8));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_yt_rsc_0_0_cgo_cse <= '0';
        reg_yt_rsc_0_16_cgo_cse <= '0';
        reg_yt_rsc_1_0_cgo_cse <= '0';
        reg_yt_rsc_1_16_cgo_cse <= '0';
        reg_xt_rsc_0_0_i_oswt_cse <= '0';
        reg_xt_rsc_0_16_i_oswt_cse <= '0';
        reg_xt_rsc_1_0_i_oswt_cse <= '0';
        reg_xt_rsc_1_16_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_0_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_1_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_2_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_3_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_4_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_5_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_6_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_7_i_oswt_cse <= '0';
        reg_twiddle_rsc_0_8_i_oswt_cse <= '0';
        twiddle_h_rsc_0_0_i_s_raddr_core_4 <= '0';
        reg_xt_rsc_triosy_1_31_obj_iswt0_cse <= '0';
        reg_ensig_cgo_cse <= '0';
        reg_ensig_cgo_17_cse <= '0';
        butterFly2_19_tw_asn_itm <= STD_LOGIC_VECTOR'( "00");
        INNER_LOOP1_stage_0 <= '0';
        INNER_LOOP1_r_9_4_sva_4_0 <= STD_LOGIC_VECTOR'( "00000");
        INNER_LOOP1_stage_0_2 <= '0';
        INNER_LOOP1_stage_0_3 <= '0';
        INNER_LOOP1_stage_0_4 <= '0';
        INNER_LOOP1_stage_0_5 <= '0';
        INNER_LOOP1_stage_0_6 <= '0';
        INNER_LOOP1_stage_0_7 <= '0';
        INNER_LOOP1_stage_0_8 <= '0';
        INNER_LOOP1_stage_0_9 <= '0';
        INNER_LOOP1_stage_0_10 <= '0';
        INNER_LOOP1_stage_0_11 <= '0';
        INNER_LOOP1_stage_0_12 <= '0';
        INNER_LOOP1_stage_0_13 <= '0';
        INNER_LOOP2_stage_0 <= '0';
        INNER_LOOP2_r_9_4_sva_4_0 <= STD_LOGIC_VECTOR'( "00000");
        INNER_LOOP2_stage_0_2 <= '0';
        INNER_LOOP2_stage_0_3 <= '0';
        INNER_LOOP2_stage_0_4 <= '0';
        INNER_LOOP2_stage_0_5 <= '0';
        INNER_LOOP2_stage_0_6 <= '0';
        INNER_LOOP2_stage_0_7 <= '0';
        INNER_LOOP2_stage_0_8 <= '0';
        INNER_LOOP2_stage_0_9 <= '0';
        INNER_LOOP2_stage_0_10 <= '0';
        INNER_LOOP2_stage_0_11 <= '0';
        INNER_LOOP2_stage_0_12 <= '0';
        INNER_LOOP3_stage_0 <= '0';
        INNER_LOOP3_r_9_4_sva_4_0 <= STD_LOGIC_VECTOR'( "00000");
        INNER_LOOP3_stage_0_2 <= '0';
        INNER_LOOP3_stage_0_3 <= '0';
        INNER_LOOP3_stage_0_4 <= '0';
        INNER_LOOP3_stage_0_5 <= '0';
        INNER_LOOP3_stage_0_6 <= '0';
        INNER_LOOP3_stage_0_7 <= '0';
        INNER_LOOP3_stage_0_8 <= '0';
        INNER_LOOP3_stage_0_9 <= '0';
        INNER_LOOP3_stage_0_10 <= '0';
        INNER_LOOP3_stage_0_11 <= '0';
        INNER_LOOP3_stage_0_12 <= '0';
        INNER_LOOP3_stage_0_13 <= '0';
        INNER_LOOP4_stage_0 <= '0';
        INNER_LOOP4_r_9_4_sva_4_0 <= STD_LOGIC_VECTOR'( "00000");
        INNER_LOOP4_stage_0_2 <= '0';
        INNER_LOOP4_stage_0_3 <= '0';
        INNER_LOOP4_stage_0_4 <= '0';
        INNER_LOOP4_stage_0_5 <= '0';
        INNER_LOOP4_stage_0_6 <= '0';
        INNER_LOOP4_stage_0_7 <= '0';
        INNER_LOOP4_stage_0_8 <= '0';
        INNER_LOOP4_stage_0_9 <= '0';
        INNER_LOOP4_stage_0_10 <= '0';
        INNER_LOOP4_stage_0_11 <= '0';
        INNER_LOOP4_stage_0_12 <= '0';
      ELSIF ( core_wen = '1' ) THEN
        reg_yt_rsc_0_0_cgo_cse <= or_67_rmff;
        reg_yt_rsc_0_16_cgo_cse <= or_166_rmff;
        reg_yt_rsc_1_0_cgo_cse <= or_248_rmff;
        reg_yt_rsc_1_16_cgo_cse <= or_347_rmff;
        reg_xt_rsc_0_0_i_oswt_cse <= or_429_rmff;
        reg_xt_rsc_0_16_i_oswt_cse <= or_512_rmff;
        reg_xt_rsc_1_0_i_oswt_cse <= or_578_rmff;
        reg_xt_rsc_1_16_i_oswt_cse <= or_660_rmff;
        reg_twiddle_rsc_0_0_i_oswt_cse <= INNER_LOOP3_INNER_LOOP3_and_1_cse OR and_1665_cse
            OR and_1666_cse OR INNER_LOOP4_INNER_LOOP4_and_1_cse;
        reg_twiddle_rsc_0_1_i_oswt_cse <= (and_dcpl_174 AND (fsm_output(6))) OR and_1686_cse;
        reg_twiddle_rsc_0_2_i_oswt_cse <= (and_dcpl_176 AND (fsm_output(6))) OR and_1695_cse;
        reg_twiddle_rsc_0_3_i_oswt_cse <= (and_dcpl_174 AND (operator_33_true_2_lshift_psp_2_0_sva(1))
            AND (fsm_output(6))) OR and_1704_cse;
        reg_twiddle_rsc_0_4_i_oswt_cse <= (INNER_LOOP3_stage_0 AND (operator_33_true_2_lshift_psp_2_0_sva(2))
            AND (fsm_output(6))) OR INNER_LOOP4_INNER_LOOP4_and_1_cse;
        reg_twiddle_rsc_0_5_i_oswt_cse <= (and_dcpl_174 AND (operator_33_true_2_lshift_psp_2_0_sva(2))
            AND (fsm_output(6))) OR and_1686_cse;
        reg_twiddle_rsc_0_6_i_oswt_cse <= (and_dcpl_176 AND (operator_33_true_2_lshift_psp_2_0_sva(2))
            AND (fsm_output(6))) OR and_1695_cse;
        reg_twiddle_rsc_0_7_i_oswt_cse <= (and_dcpl_174 AND CONV_SL_1_1(operator_33_true_2_lshift_psp_2_0_sva(2
            DOWNTO 1)=STD_LOGIC_VECTOR'("11")) AND (fsm_output(6))) OR and_1704_cse;
        reg_twiddle_rsc_0_8_i_oswt_cse <= INNER_LOOP3_INNER_LOOP3_and_1_cse OR INNER_LOOP4_INNER_LOOP4_and_1_cse;
        twiddle_h_rsc_0_0_i_s_raddr_core_4 <= MUX1HOT_s_1_4_2((INNER_LOOP1_tw_and_psp_sva_1(4)),
            (INNER_LOOP2_r_9_4_sva_4_0(4)), (INNER_LOOP3_r_9_4_sva_4_0(4)), (INNER_LOOP4_r_9_4_sva_4_0(4)),
            STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6))
            & (fsm_output(8))));
        reg_xt_rsc_triosy_1_31_obj_iswt0_cse <= and_dcpl_144 AND (fsm_output(8));
        reg_ensig_cgo_cse <= or_833_rmff;
        reg_ensig_cgo_17_cse <= or_956_rmff;
        butterFly2_19_tw_asn_itm <= MUX1HOT_v_2_4_2(STD_LOGIC_VECTOR'( "10"), (operator_20_false_acc_cse_sva(2
            DOWNTO 1)), operator_33_true_3_lshift_psp_1_0_sva_mx0w2, operator_33_true_3_lshift_psp_1_0_sva,
            STD_LOGIC_VECTOR'( nor_4_nl & (fsm_output(4)) & (fsm_output(7)) & (fsm_output(8))));
        INNER_LOOP1_stage_0 <= NOT((NOT(INNER_LOOP1_stage_0 AND (NOT (INNER_LOOP1_r_9_4_sva_2(5)))))
            AND (fsm_output(2)));
        INNER_LOOP1_r_9_4_sva_4_0 <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), (INNER_LOOP1_r_9_4_sva_2(4
            DOWNTO 0)), (fsm_output(2)));
        INNER_LOOP1_stage_0_2 <= and_1665_cse;
        INNER_LOOP1_stage_0_3 <= INNER_LOOP1_stage_0_2 AND (fsm_output(2));
        INNER_LOOP1_stage_0_4 <= INNER_LOOP1_stage_0_3 AND (fsm_output(2));
        INNER_LOOP1_stage_0_5 <= INNER_LOOP1_stage_0_4 AND (fsm_output(2));
        INNER_LOOP1_stage_0_6 <= INNER_LOOP1_stage_0_5 AND (fsm_output(2));
        INNER_LOOP1_stage_0_7 <= INNER_LOOP1_stage_0_6 AND (fsm_output(2));
        INNER_LOOP1_stage_0_8 <= INNER_LOOP1_stage_0_7 AND (fsm_output(2));
        INNER_LOOP1_stage_0_9 <= INNER_LOOP1_stage_0_8 AND (fsm_output(2));
        INNER_LOOP1_stage_0_10 <= INNER_LOOP1_stage_0_9 AND (fsm_output(2));
        INNER_LOOP1_stage_0_11 <= INNER_LOOP1_stage_0_10 AND (fsm_output(2));
        INNER_LOOP1_stage_0_12 <= INNER_LOOP1_stage_0_11 AND (fsm_output(2));
        INNER_LOOP1_stage_0_13 <= INNER_LOOP1_stage_0_12 AND (fsm_output(2));
        INNER_LOOP2_stage_0 <= NOT((NOT(INNER_LOOP2_stage_0 AND (NOT (z_out_33(5)))))
            AND (fsm_output(4)));
        INNER_LOOP2_r_9_4_sva_4_0 <= INNER_LOOP1_r_INNER_LOOP1_r_and_2_cse;
        INNER_LOOP2_stage_0_2 <= and_1666_cse;
        INNER_LOOP2_stage_0_3 <= INNER_LOOP2_stage_0_2 AND (fsm_output(4));
        INNER_LOOP2_stage_0_4 <= INNER_LOOP2_stage_0_3 AND (fsm_output(4));
        INNER_LOOP2_stage_0_5 <= INNER_LOOP2_stage_0_4 AND (fsm_output(4));
        INNER_LOOP2_stage_0_6 <= INNER_LOOP2_stage_0_5 AND (fsm_output(4));
        INNER_LOOP2_stage_0_7 <= INNER_LOOP2_stage_0_6 AND (fsm_output(4));
        INNER_LOOP2_stage_0_8 <= INNER_LOOP2_stage_0_7 AND (fsm_output(4));
        INNER_LOOP2_stage_0_9 <= INNER_LOOP2_stage_0_8 AND (fsm_output(4));
        INNER_LOOP2_stage_0_10 <= INNER_LOOP2_stage_0_9 AND (fsm_output(4));
        INNER_LOOP2_stage_0_11 <= INNER_LOOP2_stage_0_10 AND (fsm_output(4));
        INNER_LOOP2_stage_0_12 <= INNER_LOOP2_stage_0_11 AND (fsm_output(4));
        INNER_LOOP3_stage_0 <= NOT((NOT(INNER_LOOP3_stage_0 AND (NOT (z_out_33(5)))))
            AND (fsm_output(6)));
        INNER_LOOP3_r_9_4_sva_4_0 <= MUX_v_5_2_2(STD_LOGIC_VECTOR'("00000"), (z_out_33(4
            DOWNTO 0)), (fsm_output(6)));
        INNER_LOOP3_stage_0_2 <= INNER_LOOP3_INNER_LOOP3_and_1_cse;
        INNER_LOOP3_stage_0_3 <= INNER_LOOP3_stage_0_2 AND (fsm_output(6));
        INNER_LOOP3_stage_0_4 <= INNER_LOOP3_stage_0_3 AND (fsm_output(6));
        INNER_LOOP3_stage_0_5 <= INNER_LOOP3_stage_0_4 AND (fsm_output(6));
        INNER_LOOP3_stage_0_6 <= INNER_LOOP3_stage_0_5 AND (fsm_output(6));
        INNER_LOOP3_stage_0_7 <= INNER_LOOP3_stage_0_6 AND (fsm_output(6));
        INNER_LOOP3_stage_0_8 <= INNER_LOOP3_stage_0_7 AND (fsm_output(6));
        INNER_LOOP3_stage_0_9 <= INNER_LOOP3_stage_0_8 AND (fsm_output(6));
        INNER_LOOP3_stage_0_10 <= INNER_LOOP3_stage_0_9 AND (fsm_output(6));
        INNER_LOOP3_stage_0_11 <= INNER_LOOP3_stage_0_10 AND (fsm_output(6));
        INNER_LOOP3_stage_0_12 <= INNER_LOOP3_stage_0_11 AND (fsm_output(6));
        INNER_LOOP3_stage_0_13 <= INNER_LOOP3_stage_0_12 AND (fsm_output(6));
        INNER_LOOP4_stage_0 <= NOT((NOT(INNER_LOOP4_stage_0 AND (NOT (INNER_LOOP4_r_9_4_sva_2(5)))))
            AND (fsm_output(8)));
        INNER_LOOP4_r_9_4_sva_4_0 <= INNER_LOOP1_r_INNER_LOOP1_r_and_6_cse;
        INNER_LOOP4_stage_0_2 <= INNER_LOOP4_INNER_LOOP4_and_1_cse;
        INNER_LOOP4_stage_0_3 <= INNER_LOOP4_stage_0_2 AND (fsm_output(8));
        INNER_LOOP4_stage_0_4 <= INNER_LOOP4_stage_0_3 AND (fsm_output(8));
        INNER_LOOP4_stage_0_5 <= INNER_LOOP4_stage_0_4 AND (fsm_output(8));
        INNER_LOOP4_stage_0_6 <= INNER_LOOP4_stage_0_5 AND (fsm_output(8));
        INNER_LOOP4_stage_0_7 <= INNER_LOOP4_stage_0_6 AND (fsm_output(8));
        INNER_LOOP4_stage_0_8 <= INNER_LOOP4_stage_0_7 AND (fsm_output(8));
        INNER_LOOP4_stage_0_9 <= INNER_LOOP4_stage_0_8 AND (fsm_output(8));
        INNER_LOOP4_stage_0_10 <= INNER_LOOP4_stage_0_9 AND (fsm_output(8));
        INNER_LOOP4_stage_0_11 <= INNER_LOOP4_stage_0_10 AND (fsm_output(8));
        INNER_LOOP4_stage_0_12 <= INNER_LOOP4_stage_0_11 AND (fsm_output(8));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_160_itm_12 <= '0';
      ELSIF ( (core_wen AND INNER_LOOP1_stage_0_12) = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_160_itm_12 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_11;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( modulo_add_qelse_and_cse = '1' ) THEN
        modulo_add_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_sva_1, z_out_87,
            z_out_32_1);
        modulo_add_1_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_1_sva_1, z_out_88,
            z_out_1_32);
        modulo_add_2_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_2_sva_1, z_out_89,
            z_out_2_32);
        modulo_add_3_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_3_sva_1, z_out_90,
            z_out_3_32);
        modulo_add_4_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_4_sva_1, z_out_91,
            z_out_4_32);
        modulo_add_5_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_5_sva_1, z_out_92,
            z_out_5_32);
        modulo_add_6_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_6_sva_1, z_out_93,
            z_out_6_32);
        modulo_add_7_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_7_sva_1, z_out_94,
            z_out_7_32);
        modulo_add_8_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_8_sva_1, z_out_95,
            z_out_8_32);
        modulo_add_9_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_9_sva_1, z_out_96,
            z_out_9_32);
        modulo_add_10_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_10_sva_1, z_out_97,
            z_out_10_32);
        modulo_add_11_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_11_sva_1, z_out_98,
            z_out_11_32);
        modulo_add_12_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_12_sva_1, z_out_99,
            z_out_12_32);
        modulo_add_13_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_13_sva_1, z_out_100,
            z_out_13_32);
        modulo_add_14_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_14_sva_1, z_out_101,
            z_out_14_32);
        modulo_add_15_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_15_sva_1, z_out_102,
            z_out_15_32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_11 <= '0';
      ELSIF ( modulo_add_qelse_and_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_11 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_10;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_11 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_10))
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_290_itm_11 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_385_itm_10;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_11 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_10)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_306_itm_11 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_401_itm_10;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly1_and_cse = '1' ) THEN
        modulo_add_base_15_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_94_lpi_3_dfm_8)
            + UNSIGNED(mult_15_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_14_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_92_lpi_3_dfm_8)
            + UNSIGNED(mult_14_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_13_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_90_lpi_3_dfm_8)
            + UNSIGNED(mult_13_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_12_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_88_lpi_3_dfm_8)
            + UNSIGNED(mult_12_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_11_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_86_lpi_3_dfm_8)
            + UNSIGNED(mult_11_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_10_sva_1 <= z_out_85;
        modulo_add_base_9_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_82_lpi_3_dfm_8)
            + UNSIGNED(mult_9_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_8_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_80_lpi_3_dfm_8)
            + UNSIGNED(mult_8_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_7_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_78_lpi_3_dfm_8)
            + UNSIGNED(mult_7_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_6_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_76_lpi_3_dfm_8)
            + UNSIGNED(mult_6_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_5_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_74_lpi_3_dfm_8)
            + UNSIGNED(mult_5_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_4_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_72_lpi_3_dfm_8)
            + UNSIGNED(mult_4_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_3_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_70_lpi_3_dfm_8)
            + UNSIGNED(mult_3_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_2_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_68_lpi_3_dfm_8)
            + UNSIGNED(mult_2_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_1_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_66_lpi_3_dfm_8)
            + UNSIGNED(mult_1_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_64_lpi_3_dfm_8)
            + UNSIGNED(mult_res_lpi_3_dfm_mx0), 32));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        modulo_sub_base_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_1_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_2_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_3_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_4_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_5_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_6_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_7_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_8_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_9_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_10_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_11_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_12_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_13_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_14_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_15_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_10 <= '0';
      ELSIF ( butterFly1_and_cse = '1' ) THEN
        modulo_sub_base_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_64_lpi_3_dfm_8)
            - SIGNED(mult_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_1_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_66_lpi_3_dfm_8)
            - SIGNED(mult_1_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_2_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_68_lpi_3_dfm_8)
            - SIGNED(mult_2_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_3_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_70_lpi_3_dfm_8)
            - SIGNED(mult_3_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_4_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_72_lpi_3_dfm_8)
            - SIGNED(mult_4_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_5_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_74_lpi_3_dfm_8)
            - SIGNED(mult_5_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_6_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_76_lpi_3_dfm_8)
            - SIGNED(mult_6_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_7_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_78_lpi_3_dfm_8)
            - SIGNED(mult_7_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_8_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_80_lpi_3_dfm_8)
            - SIGNED(mult_8_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_9_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_82_lpi_3_dfm_8)
            - SIGNED(mult_9_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_10_sva_1 <= z_out_86;
        modulo_sub_base_11_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_86_lpi_3_dfm_8)
            - SIGNED(mult_11_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_12_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_88_lpi_3_dfm_8)
            - SIGNED(mult_12_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_13_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_90_lpi_3_dfm_8)
            - SIGNED(mult_13_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_14_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_92_lpi_3_dfm_8)
            - SIGNED(mult_14_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_15_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_94_lpi_3_dfm_8)
            - SIGNED(mult_15_res_lpi_3_dfm_mx0), 32));
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_10 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_10 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_9))
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_385_itm_10 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_10 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_9)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_401_itm_10 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_15_if_and_cse = '1' ) THEN
        mult_res_sva_1 <= mult_res_sva_2;
        mult_1_res_sva_1 <= mult_1_res_sva_2;
        mult_2_res_sva_1 <= mult_2_res_sva_2;
        mult_3_res_sva_1 <= mult_3_res_sva_2;
        mult_4_res_sva_1 <= mult_4_res_sva_2;
        mult_5_res_sva_1 <= mult_5_res_sva_2;
        mult_6_res_sva_1 <= mult_6_res_sva_2;
        mult_7_res_sva_1 <= mult_7_res_sva_2;
        mult_8_res_sva_1 <= mult_8_res_sva_2;
        mult_9_res_sva_1 <= mult_9_res_sva_2;
        mult_10_res_sva_1 <= mult_10_res_sva_2;
        mult_11_res_sva_1 <= mult_11_res_sva_2;
        mult_12_res_sva_1 <= mult_12_res_sva_2;
        mult_13_res_sva_1 <= mult_13_res_sva_2;
        mult_14_res_sva_1 <= mult_14_res_sva_2;
        mult_15_res_sva_1 <= mult_15_res_sva_2;
        tmp_94_lpi_3_dfm_8 <= tmp_94_lpi_3_dfm_7;
        tmp_92_lpi_3_dfm_8 <= tmp_92_lpi_3_dfm_7;
        tmp_90_lpi_3_dfm_8 <= tmp_90_lpi_3_dfm_7;
        tmp_88_lpi_3_dfm_8 <= tmp_88_lpi_3_dfm_7;
        tmp_86_lpi_3_dfm_8 <= tmp_86_lpi_3_dfm_7;
        tmp_84_lpi_3_dfm_8 <= tmp_84_lpi_3_dfm_7;
        tmp_82_lpi_3_dfm_8 <= tmp_82_lpi_3_dfm_7;
        tmp_80_lpi_3_dfm_8 <= tmp_80_lpi_3_dfm_7;
        tmp_78_lpi_3_dfm_8 <= tmp_78_lpi_3_dfm_7;
        tmp_76_lpi_3_dfm_8 <= tmp_76_lpi_3_dfm_7;
        tmp_74_lpi_3_dfm_8 <= tmp_74_lpi_3_dfm_7;
        tmp_72_lpi_3_dfm_8 <= tmp_72_lpi_3_dfm_7;
        tmp_70_lpi_3_dfm_8 <= tmp_70_lpi_3_dfm_7;
        tmp_68_lpi_3_dfm_8 <= tmp_68_lpi_3_dfm_7;
        tmp_66_lpi_3_dfm_8 <= tmp_66_lpi_3_dfm_7;
        tmp_64_lpi_3_dfm_8 <= tmp_64_lpi_3_dfm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        mult_15_slc_32_svs_st_1 <= '0';
        mult_14_slc_32_svs_st_1 <= '0';
        mult_13_slc_32_svs_st_1 <= '0';
        mult_12_slc_32_svs_st_1 <= '0';
        mult_11_slc_32_svs_st_1 <= '0';
        mult_10_slc_32_svs_st_1 <= '0';
        mult_9_slc_32_svs_st_1 <= '0';
        mult_8_slc_32_svs_st_1 <= '0';
        mult_7_slc_32_svs_st_1 <= '0';
        mult_6_slc_32_svs_st_1 <= '0';
        mult_5_slc_32_svs_st_1 <= '0';
        mult_4_slc_32_svs_st_1 <= '0';
        mult_3_slc_32_svs_st_1 <= '0';
        mult_2_slc_32_svs_st_1 <= '0';
        mult_1_slc_32_svs_st_1 <= '0';
        mult_slc_32_svs_st_1 <= '0';
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_9 <= '0';
      ELSIF ( mult_15_if_and_cse = '1' ) THEN
        mult_15_slc_32_svs_st_1 <= z_out_16_32;
        mult_14_slc_32_svs_st_1 <= z_out_17_32;
        mult_13_slc_32_svs_st_1 <= z_out_18_32;
        mult_12_slc_32_svs_st_1 <= z_out_19_32;
        mult_11_slc_32_svs_st_1 <= z_out_20_32;
        mult_10_slc_32_svs_st_1 <= z_out_21_32;
        mult_9_slc_32_svs_st_1 <= z_out_22_32;
        mult_8_slc_32_svs_st_1 <= z_out_23_32;
        mult_7_slc_32_svs_st_1 <= z_out_24_32;
        mult_6_slc_32_svs_st_1 <= z_out_25_32;
        mult_5_slc_32_svs_st_1 <= z_out_26_32;
        mult_4_slc_32_svs_st_1 <= z_out_27_32;
        mult_3_slc_32_svs_st_1 <= z_out_28_32;
        mult_2_slc_32_svs_st_1 <= z_out_29_32;
        mult_1_slc_32_svs_st_1 <= z_out_30_32;
        mult_slc_32_svs_st_1 <= z_out_31_32;
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_9 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1 <= '0';
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_1 <= '0';
      ELSIF ( INNER_LOOP1_r_and_7_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1 <= INNER_LOOP1_r_9_4_sva_4_0(4);
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_1 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND (NOT (fsm_output(2)))) = '1' ) THEN
        operator_33_true_return_8_4_sva <= z_out_32(8 DOWNTO 4);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_20_false_acc_cse_sva <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( (core_wen AND CONV_SL_1_1(fsm_output(4 DOWNTO 2)=STD_LOGIC_VECTOR'("000")))
          = '1' ) THEN
        operator_20_false_acc_cse_sva <= operator_20_false_acc_cse_sva_mx0w0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_15_z_and_cse = '1' ) THEN
        mult_15_z_asn_itm_4 <= mult_15_z_asn_itm_3;
        mult_14_z_asn_itm_4 <= mult_14_z_asn_itm_3;
        mult_13_z_asn_itm_4 <= mult_13_z_asn_itm_3;
        mult_12_z_asn_itm_4 <= mult_12_z_asn_itm_3;
        mult_11_z_asn_itm_4 <= mult_11_z_asn_itm_3;
        mult_10_z_asn_itm_4 <= mult_10_z_asn_itm_3;
        mult_9_z_asn_itm_4 <= mult_9_z_asn_itm_3;
        mult_8_z_asn_itm_4 <= mult_8_z_asn_itm_3;
        mult_7_z_asn_itm_4 <= mult_7_z_asn_itm_3;
        mult_6_z_asn_itm_4 <= mult_6_z_asn_itm_3;
        mult_5_z_asn_itm_4 <= mult_5_z_asn_itm_3;
        mult_4_z_asn_itm_4 <= mult_4_z_asn_itm_3;
        mult_3_z_asn_itm_4 <= mult_3_z_asn_itm_3;
        mult_2_z_asn_itm_4 <= mult_2_z_asn_itm_3;
        mult_1_z_asn_itm_4 <= mult_1_z_asn_itm_3;
        mult_z_asn_itm_4 <= mult_z_asn_itm_3;
        tmp_94_lpi_3_dfm_7 <= tmp_94_lpi_3_dfm_6;
        tmp_92_lpi_3_dfm_7 <= tmp_92_lpi_3_dfm_6;
        tmp_90_lpi_3_dfm_7 <= tmp_90_lpi_3_dfm_6;
        tmp_88_lpi_3_dfm_7 <= tmp_88_lpi_3_dfm_6;
        tmp_86_lpi_3_dfm_7 <= tmp_86_lpi_3_dfm_6;
        tmp_84_lpi_3_dfm_7 <= tmp_84_lpi_3_dfm_6;
        tmp_82_lpi_3_dfm_7 <= tmp_82_lpi_3_dfm_6;
        tmp_80_lpi_3_dfm_7 <= tmp_80_lpi_3_dfm_6;
        tmp_78_lpi_3_dfm_7 <= tmp_78_lpi_3_dfm_6;
        tmp_76_lpi_3_dfm_7 <= tmp_76_lpi_3_dfm_6;
        tmp_74_lpi_3_dfm_7 <= tmp_74_lpi_3_dfm_6;
        tmp_72_lpi_3_dfm_7 <= tmp_72_lpi_3_dfm_6;
        tmp_70_lpi_3_dfm_7 <= tmp_70_lpi_3_dfm_6;
        tmp_68_lpi_3_dfm_7 <= tmp_68_lpi_3_dfm_6;
        tmp_66_lpi_3_dfm_7 <= tmp_66_lpi_3_dfm_6;
        tmp_64_lpi_3_dfm_7 <= tmp_64_lpi_3_dfm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_8 <= '0';
      ELSIF ( mult_15_z_and_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_15_z_and_cse_1 = '1' ) THEN
        reg_mult_15_z_asn_itm_1_cse <= mult_z_mul_cmp_1_z;
        reg_mult_14_z_asn_itm_1_cse <= mult_z_mul_cmp_3_z;
        reg_mult_13_z_asn_itm_1_cse <= mult_z_mul_cmp_5_z;
        reg_mult_12_z_asn_itm_1_cse <= mult_z_mul_cmp_7_z;
        reg_mult_11_z_asn_itm_1_cse <= mult_z_mul_cmp_9_z;
        reg_mult_10_z_asn_itm_1_cse <= mult_z_mul_cmp_11_z;
        reg_mult_9_z_asn_itm_1_cse <= mult_z_mul_cmp_13_z;
        reg_mult_8_z_asn_itm_1_cse <= mult_z_mul_cmp_15_z;
        reg_mult_7_z_asn_itm_1_cse <= mult_z_mul_cmp_17_z;
        reg_mult_6_z_asn_itm_1_cse <= mult_z_mul_cmp_19_z;
        reg_mult_5_z_asn_itm_1_cse <= mult_z_mul_cmp_21_z;
        reg_mult_4_z_asn_itm_1_cse <= mult_z_mul_cmp_23_z;
        reg_mult_3_z_asn_itm_1_cse <= mult_z_mul_cmp_25_z;
        reg_mult_2_z_asn_itm_1_cse <= mult_z_mul_cmp_27_z;
        reg_mult_1_z_asn_itm_1_cse <= mult_z_mul_cmp_29_z;
        reg_mult_z_asn_itm_1_cse <= mult_z_mul_cmp_31_z;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_9 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_8)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_9 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_9 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_8))
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_9 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_8 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_7)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_8 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_7))
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_8 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_15_z_and_1_cse = '1' ) THEN
        mult_15_z_asn_itm_3 <= mult_15_z_asn_itm_2;
        mult_14_z_asn_itm_3 <= mult_14_z_asn_itm_2;
        mult_13_z_asn_itm_3 <= mult_13_z_asn_itm_2;
        mult_12_z_asn_itm_3 <= mult_12_z_asn_itm_2;
        mult_11_z_asn_itm_3 <= mult_11_z_asn_itm_2;
        mult_10_z_asn_itm_3 <= mult_10_z_asn_itm_2;
        mult_9_z_asn_itm_3 <= mult_9_z_asn_itm_2;
        mult_8_z_asn_itm_3 <= mult_8_z_asn_itm_2;
        mult_7_z_asn_itm_3 <= mult_7_z_asn_itm_2;
        mult_6_z_asn_itm_3 <= mult_6_z_asn_itm_2;
        mult_5_z_asn_itm_3 <= mult_5_z_asn_itm_2;
        mult_4_z_asn_itm_3 <= mult_4_z_asn_itm_2;
        mult_3_z_asn_itm_3 <= mult_3_z_asn_itm_2;
        mult_2_z_asn_itm_3 <= mult_2_z_asn_itm_2;
        mult_1_z_asn_itm_3 <= mult_1_z_asn_itm_2;
        mult_z_asn_itm_3 <= mult_z_asn_itm_2;
        tmp_94_lpi_3_dfm_6 <= tmp_94_lpi_3_dfm_5;
        tmp_92_lpi_3_dfm_6 <= tmp_92_lpi_3_dfm_5;
        tmp_90_lpi_3_dfm_6 <= tmp_90_lpi_3_dfm_5;
        tmp_88_lpi_3_dfm_6 <= tmp_88_lpi_3_dfm_5;
        tmp_86_lpi_3_dfm_6 <= tmp_86_lpi_3_dfm_5;
        tmp_84_lpi_3_dfm_6 <= tmp_84_lpi_3_dfm_5;
        tmp_82_lpi_3_dfm_6 <= tmp_82_lpi_3_dfm_5;
        tmp_80_lpi_3_dfm_6 <= tmp_80_lpi_3_dfm_5;
        tmp_78_lpi_3_dfm_6 <= tmp_78_lpi_3_dfm_5;
        tmp_76_lpi_3_dfm_6 <= tmp_76_lpi_3_dfm_5;
        tmp_74_lpi_3_dfm_6 <= tmp_74_lpi_3_dfm_5;
        tmp_72_lpi_3_dfm_6 <= tmp_72_lpi_3_dfm_5;
        tmp_70_lpi_3_dfm_6 <= tmp_70_lpi_3_dfm_5;
        tmp_68_lpi_3_dfm_6 <= tmp_68_lpi_3_dfm_5;
        tmp_66_lpi_3_dfm_6 <= tmp_66_lpi_3_dfm_5;
        tmp_64_lpi_3_dfm_6 <= tmp_64_lpi_3_dfm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_7 <= '0';
      ELSIF ( mult_15_z_and_1_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_7 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_6)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_7 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_6))
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_7 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_15_z_and_2_cse = '1' ) THEN
        mult_15_z_asn_itm_2 <= mult_15_z_asn_itm_1;
        mult_14_z_asn_itm_2 <= mult_14_z_asn_itm_1;
        mult_13_z_asn_itm_2 <= mult_13_z_asn_itm_1;
        mult_12_z_asn_itm_2 <= mult_12_z_asn_itm_1;
        mult_11_z_asn_itm_2 <= mult_11_z_asn_itm_1;
        mult_10_z_asn_itm_2 <= mult_10_z_asn_itm_1;
        mult_9_z_asn_itm_2 <= mult_9_z_asn_itm_1;
        mult_8_z_asn_itm_2 <= mult_8_z_asn_itm_1;
        mult_7_z_asn_itm_2 <= mult_7_z_asn_itm_1;
        mult_6_z_asn_itm_2 <= mult_6_z_asn_itm_1;
        mult_5_z_asn_itm_2 <= mult_5_z_asn_itm_1;
        mult_4_z_asn_itm_2 <= mult_4_z_asn_itm_1;
        mult_3_z_asn_itm_2 <= mult_3_z_asn_itm_1;
        mult_2_z_asn_itm_2 <= mult_2_z_asn_itm_1;
        mult_1_z_asn_itm_2 <= mult_1_z_asn_itm_1;
        mult_z_asn_itm_2 <= mult_z_asn_itm_1;
        tmp_94_lpi_3_dfm_5 <= tmp_94_lpi_3_dfm_4;
        tmp_92_lpi_3_dfm_5 <= tmp_92_lpi_3_dfm_4;
        tmp_90_lpi_3_dfm_5 <= tmp_90_lpi_3_dfm_4;
        tmp_88_lpi_3_dfm_5 <= tmp_88_lpi_3_dfm_4;
        tmp_86_lpi_3_dfm_5 <= tmp_86_lpi_3_dfm_4;
        tmp_84_lpi_3_dfm_5 <= tmp_84_lpi_3_dfm_4;
        tmp_82_lpi_3_dfm_5 <= tmp_82_lpi_3_dfm_4;
        tmp_80_lpi_3_dfm_5 <= tmp_80_lpi_3_dfm_4;
        tmp_78_lpi_3_dfm_5 <= tmp_78_lpi_3_dfm_4;
        tmp_76_lpi_3_dfm_5 <= tmp_76_lpi_3_dfm_4;
        tmp_74_lpi_3_dfm_5 <= tmp_74_lpi_3_dfm_4;
        tmp_72_lpi_3_dfm_5 <= tmp_72_lpi_3_dfm_4;
        tmp_70_lpi_3_dfm_5 <= tmp_70_lpi_3_dfm_4;
        tmp_68_lpi_3_dfm_5 <= tmp_68_lpi_3_dfm_4;
        tmp_66_lpi_3_dfm_5 <= tmp_66_lpi_3_dfm_4;
        tmp_64_lpi_3_dfm_5 <= tmp_64_lpi_3_dfm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_6 <= '0';
      ELSIF ( mult_15_z_and_2_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_6 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_5)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_6 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_5))
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_6 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_15_z_and_3_cse = '1' ) THEN
        mult_15_z_asn_itm_1 <= mult_z_mul_cmp_2_z;
        mult_14_z_asn_itm_1 <= mult_z_mul_cmp_4_z;
        mult_13_z_asn_itm_1 <= mult_z_mul_cmp_6_z;
        mult_12_z_asn_itm_1 <= mult_z_mul_cmp_8_z;
        mult_11_z_asn_itm_1 <= mult_z_mul_cmp_10_z;
        mult_10_z_asn_itm_1 <= mult_z_mul_cmp_12_z;
        mult_9_z_asn_itm_1 <= mult_z_mul_cmp_14_z;
        mult_8_z_asn_itm_1 <= mult_z_mul_cmp_16_z;
        mult_7_z_asn_itm_1 <= mult_z_mul_cmp_18_z;
        mult_6_z_asn_itm_1 <= mult_z_mul_cmp_20_z;
        mult_5_z_asn_itm_1 <= mult_z_mul_cmp_22_z;
        mult_4_z_asn_itm_1 <= mult_z_mul_cmp_24_z;
        mult_3_z_asn_itm_1 <= mult_z_mul_cmp_26_z;
        mult_2_z_asn_itm_1 <= mult_z_mul_cmp_28_z;
        mult_1_z_asn_itm_1 <= mult_z_mul_cmp_30_z;
        mult_z_asn_itm_1 <= mult_z_mul_cmp_z;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP1_r_and_20_cse = '1' ) THEN
        tmp_94_lpi_3_dfm_4 <= tmp_94_lpi_3_dfm_3;
        tmp_92_lpi_3_dfm_4 <= tmp_92_lpi_3_dfm_3;
        tmp_90_lpi_3_dfm_4 <= tmp_90_lpi_3_dfm_3;
        tmp_88_lpi_3_dfm_4 <= tmp_88_lpi_3_dfm_3;
        tmp_86_lpi_3_dfm_4 <= tmp_86_lpi_3_dfm_3;
        tmp_84_lpi_3_dfm_4 <= tmp_84_lpi_3_dfm_3;
        tmp_82_lpi_3_dfm_4 <= tmp_82_lpi_3_dfm_3;
        tmp_80_lpi_3_dfm_4 <= tmp_80_lpi_3_dfm_3;
        tmp_78_lpi_3_dfm_4 <= tmp_78_lpi_3_dfm_3;
        tmp_76_lpi_3_dfm_4 <= tmp_76_lpi_3_dfm_3;
        tmp_74_lpi_3_dfm_4 <= tmp_74_lpi_3_dfm_3;
        tmp_72_lpi_3_dfm_4 <= tmp_72_lpi_3_dfm_3;
        tmp_70_lpi_3_dfm_4 <= tmp_70_lpi_3_dfm_3;
        tmp_68_lpi_3_dfm_4 <= tmp_68_lpi_3_dfm_3;
        tmp_66_lpi_3_dfm_4 <= tmp_66_lpi_3_dfm_3;
        tmp_64_lpi_3_dfm_4 <= tmp_64_lpi_3_dfm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_5 <= '0';
      ELSIF ( INNER_LOOP1_r_and_20_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_5 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_4)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_5 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_4))
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_5 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP1_r_and_23_cse = '1' ) THEN
        tmp_94_lpi_3_dfm_3 <= tmp_94_lpi_3_dfm_2;
        tmp_92_lpi_3_dfm_3 <= tmp_92_lpi_3_dfm_2;
        tmp_90_lpi_3_dfm_3 <= tmp_90_lpi_3_dfm_2;
        tmp_88_lpi_3_dfm_3 <= tmp_88_lpi_3_dfm_2;
        tmp_86_lpi_3_dfm_3 <= tmp_86_lpi_3_dfm_2;
        tmp_84_lpi_3_dfm_3 <= tmp_84_lpi_3_dfm_2;
        tmp_82_lpi_3_dfm_3 <= tmp_82_lpi_3_dfm_2;
        tmp_80_lpi_3_dfm_3 <= tmp_80_lpi_3_dfm_2;
        tmp_78_lpi_3_dfm_3 <= tmp_78_lpi_3_dfm_2;
        tmp_76_lpi_3_dfm_3 <= tmp_76_lpi_3_dfm_2;
        tmp_74_lpi_3_dfm_3 <= tmp_74_lpi_3_dfm_2;
        tmp_72_lpi_3_dfm_3 <= tmp_72_lpi_3_dfm_2;
        tmp_70_lpi_3_dfm_3 <= tmp_70_lpi_3_dfm_2;
        tmp_68_lpi_3_dfm_3 <= tmp_68_lpi_3_dfm_2;
        tmp_66_lpi_3_dfm_3 <= tmp_66_lpi_3_dfm_2;
        tmp_64_lpi_3_dfm_3 <= tmp_64_lpi_3_dfm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_4 <= '0';
      ELSIF ( INNER_LOOP1_r_and_23_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_4 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_3)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_4 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_3))
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_4 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP1_r_and_26_cse = '1' ) THEN
        tmp_94_lpi_3_dfm_2 <= tmp_94_lpi_3_dfm_1;
        tmp_92_lpi_3_dfm_2 <= tmp_92_lpi_3_dfm_1;
        tmp_90_lpi_3_dfm_2 <= tmp_90_lpi_3_dfm_1;
        tmp_88_lpi_3_dfm_2 <= tmp_88_lpi_3_dfm_1;
        tmp_86_lpi_3_dfm_2 <= tmp_86_lpi_3_dfm_1;
        tmp_84_lpi_3_dfm_2 <= tmp_84_lpi_3_dfm_1;
        tmp_82_lpi_3_dfm_2 <= tmp_82_lpi_3_dfm_1;
        tmp_80_lpi_3_dfm_2 <= tmp_80_lpi_3_dfm_1;
        tmp_78_lpi_3_dfm_2 <= tmp_78_lpi_3_dfm_1;
        tmp_76_lpi_3_dfm_2 <= tmp_76_lpi_3_dfm_1;
        tmp_74_lpi_3_dfm_2 <= tmp_74_lpi_3_dfm_1;
        tmp_72_lpi_3_dfm_2 <= tmp_72_lpi_3_dfm_1;
        tmp_70_lpi_3_dfm_2 <= tmp_70_lpi_3_dfm_1;
        tmp_68_lpi_3_dfm_2 <= tmp_68_lpi_3_dfm_1;
        tmp_66_lpi_3_dfm_2 <= tmp_66_lpi_3_dfm_1;
        tmp_64_lpi_3_dfm_2 <= tmp_64_lpi_3_dfm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_3 <= '0';
      ELSIF ( INNER_LOOP1_r_and_26_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_3 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_2)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_3 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_2))
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_3 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP1_r_and_29_cse = '1' ) THEN
        tmp_94_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_30_i_qa_d_mxwt, xt_rsc_1_30_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_92_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_28_i_qa_d_mxwt, xt_rsc_1_28_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_90_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_26_i_qa_d_mxwt, xt_rsc_1_26_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_88_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_24_i_qa_d_mxwt, xt_rsc_1_24_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_86_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_22_i_qa_d_mxwt, xt_rsc_1_22_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_84_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_20_i_qa_d_mxwt, xt_rsc_1_20_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_82_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_18_i_qa_d_mxwt, xt_rsc_1_18_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_80_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_16_i_qa_d_mxwt, xt_rsc_1_16_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_78_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_14_i_qa_d_mxwt, xt_rsc_1_14_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_76_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_12_i_qa_d_mxwt, xt_rsc_1_12_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_74_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_10_i_qa_d_mxwt, xt_rsc_1_10_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_72_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_8_i_qa_d_mxwt, xt_rsc_1_8_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_70_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_6_i_qa_d_mxwt, xt_rsc_1_6_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_68_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_4_i_qa_d_mxwt, xt_rsc_1_4_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_66_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_2_i_qa_d_mxwt, xt_rsc_1_2_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
        tmp_64_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_0_i_qa_d_mxwt, xt_rsc_1_0_i_qa_d_mxwt,
            INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_63_itm_1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_2 <= '0';
      ELSIF ( INNER_LOOP1_r_and_29_cse = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_2 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_1)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0_2 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm_1))
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_2 <= INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0 AND INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm)
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_20_itm_1 <= INNER_LOOP1_r_9_4_sva_4_0(4
            DOWNTO 1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP1_stage_0 AND (NOT INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm))
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_4210_itm_1 <= INNER_LOOP1_r_9_4_sva_4_0(4
            DOWNTO 1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm <= '0';
      ELSIF ( (core_wen AND ((fsm_output(1)) OR ((NOT((INNER_LOOP1_r_9_4_sva_2(5))
          OR INNER_LOOP1_nor_tmp)) AND INNER_LOOP1_stage_0 AND (fsm_output(2)))))
          = '1' ) THEN
        INNER_LOOP1_r_slc_INNER_LOOP1_r_9_4_4_0_161_itm <= (INNER_LOOP1_r_9_4_sva_2(0))
            AND (fsm_output(2));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( modulo_add_16_qelse_and_cse = '1' ) THEN
        modulo_add_16_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_16_sva_1, z_out_89,
            z_out_32_1);
        modulo_sub_16_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_16_sva_1(30
            DOWNTO 0))), z_out_50, modulo_sub_base_16_sva_1(31));
        modulo_add_17_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_17_sva_1, z_out_90,
            z_out_1_32);
        modulo_sub_17_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_17_sva_1(30
            DOWNTO 0))), z_out_52, modulo_sub_base_17_sva_1(31));
        modulo_add_18_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_18_sva_1, z_out_91,
            z_out_2_32);
        modulo_sub_18_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_18_sva_1(30
            DOWNTO 0))), z_out_54, modulo_sub_base_18_sva_1(31));
        modulo_add_19_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_19_sva_1, z_out_101,
            z_out_3_32);
        modulo_sub_19_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_19_sva_1(30
            DOWNTO 0))), z_out_56, modulo_sub_base_19_sva_1(31));
        modulo_add_20_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_20_sva_1, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_20_qif_acc_nl),
            32)), z_out_4_32);
        modulo_sub_20_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_20_sva_1(30
            DOWNTO 0))), z_out_58, modulo_sub_base_20_sva_1(31));
        modulo_add_21_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_21_sva_1, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_21_qif_acc_nl),
            32)), z_out_5_32);
        modulo_sub_21_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_21_sva_1(30
            DOWNTO 0))), z_out_60, modulo_sub_base_21_sva_1(31));
        modulo_add_22_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_22_sva_1, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_22_qif_acc_nl),
            32)), z_out_6_32);
        modulo_sub_22_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_22_sva_1(30
            DOWNTO 0))), z_out_62, modulo_sub_base_22_sva_1(31));
        modulo_add_23_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_23_sva_1, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_23_qif_acc_nl),
            32)), z_out_7_32);
        modulo_sub_23_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_23_sva_1(30
            DOWNTO 0))), z_out_64, modulo_sub_base_23_sva_1(31));
        modulo_add_24_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_24_sva_1, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_24_qif_acc_nl),
            32)), z_out_8_32);
        modulo_sub_24_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_24_sva_1(30
            DOWNTO 0))), z_out_66, modulo_sub_base_24_sva_1(31));
        modulo_add_25_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_25_sva_1, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_25_qif_acc_nl),
            32)), z_out_9_32);
        modulo_sub_25_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_25_sva_1(30
            DOWNTO 0))), z_out_68, modulo_sub_base_25_sva_1(31));
        modulo_add_26_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_26_sva_1, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_26_qif_acc_nl),
            32)), z_out_10_32);
        modulo_sub_26_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_26_sva_1(30
            DOWNTO 0))), z_out_70, modulo_sub_base_26_sva_1(31));
        modulo_add_27_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_27_sva_1, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_27_qif_acc_nl),
            32)), z_out_11_32);
        modulo_sub_27_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_27_sva_1(30
            DOWNTO 0))), z_out_72, modulo_sub_base_27_sva_1(31));
        modulo_add_28_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_28_sva_1, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_28_qif_acc_nl),
            32)), z_out_12_32);
        modulo_sub_28_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_28_sva_1(30
            DOWNTO 0))), z_out_74, modulo_sub_base_28_sva_1(31));
        modulo_add_29_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_29_sva_1, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_29_qif_acc_nl),
            32)), z_out_13_32);
        modulo_sub_29_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_29_sva_1(30
            DOWNTO 0))), z_out_76, modulo_sub_base_29_sva_1(31));
        modulo_add_30_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_30_sva_1, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_30_qif_acc_nl),
            32)), z_out_14_32);
        modulo_sub_30_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_30_sva_1(30
            DOWNTO 0))), z_out_78, modulo_sub_base_30_sva_1(31));
        modulo_add_31_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_31_sva_1, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_31_qif_acc_nl),
            32)), z_out_15_32);
        modulo_sub_31_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_31_sva_1(30
            DOWNTO 0))), z_out_80, modulo_sub_base_31_sva_1(31));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_11 <= '0';
      ELSIF ( modulo_add_16_qelse_and_cse = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_11 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_10;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_11 AND (NOT INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_10))
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_290_itm_11 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_10;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_11 AND INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_10)
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_306_itm_11 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_10;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly1_31_and_cse = '1' ) THEN
        modulo_add_base_31_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_30_lpi_3_dfm_8)
            + UNSIGNED(mult_31_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_30_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_28_lpi_3_dfm_8)
            + UNSIGNED(mult_30_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_29_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_26_lpi_3_dfm_8)
            + UNSIGNED(mult_29_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_28_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_24_lpi_3_dfm_8)
            + UNSIGNED(mult_28_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_27_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_22_lpi_3_dfm_8)
            + UNSIGNED(mult_27_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_26_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_20_lpi_3_dfm_8)
            + UNSIGNED(mult_26_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_25_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_18_lpi_3_dfm_8)
            + UNSIGNED(mult_25_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_24_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_16_lpi_3_dfm_8)
            + UNSIGNED(mult_24_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_23_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_14_lpi_3_dfm_8)
            + UNSIGNED(mult_23_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_22_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_12_lpi_3_dfm_8)
            + UNSIGNED(mult_22_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_21_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_10_lpi_3_dfm_8)
            + UNSIGNED(mult_21_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_20_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_8_lpi_3_dfm_8)
            + UNSIGNED(mult_20_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_19_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_6_lpi_3_dfm_8)
            + UNSIGNED(mult_19_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_18_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_4_lpi_3_dfm_8)
            + UNSIGNED(mult_18_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_17_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_2_lpi_3_dfm_8)
            + UNSIGNED(mult_17_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_16_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_lpi_3_dfm_8)
            + UNSIGNED(mult_16_res_lpi_3_dfm_mx0), 32));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        modulo_sub_base_16_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_17_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_18_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_19_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_20_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_21_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_22_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_23_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_24_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_25_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_26_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_27_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_28_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_29_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_30_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_31_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_10 <= '0';
      ELSIF ( butterFly1_31_and_cse = '1' ) THEN
        modulo_sub_base_16_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_lpi_3_dfm_8)
            - SIGNED(mult_16_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_17_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_2_lpi_3_dfm_8)
            - SIGNED(mult_17_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_18_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_4_lpi_3_dfm_8)
            - SIGNED(mult_18_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_19_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_6_lpi_3_dfm_8)
            - SIGNED(mult_19_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_20_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_8_lpi_3_dfm_8)
            - SIGNED(mult_20_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_21_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_10_lpi_3_dfm_8)
            - SIGNED(mult_21_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_22_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_12_lpi_3_dfm_8)
            - SIGNED(mult_22_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_23_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_14_lpi_3_dfm_8)
            - SIGNED(mult_23_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_24_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_16_lpi_3_dfm_8)
            - SIGNED(mult_24_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_25_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_18_lpi_3_dfm_8)
            - SIGNED(mult_25_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_26_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_20_lpi_3_dfm_8)
            - SIGNED(mult_26_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_27_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_22_lpi_3_dfm_8)
            - SIGNED(mult_27_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_28_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_24_lpi_3_dfm_8)
            - SIGNED(mult_28_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_29_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_26_lpi_3_dfm_8)
            - SIGNED(mult_29_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_30_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_28_lpi_3_dfm_8)
            - SIGNED(mult_30_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_31_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_30_lpi_3_dfm_8)
            - SIGNED(mult_31_res_lpi_3_dfm_mx0), 32));
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_10 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_31_if_and_cse = '1' ) THEN
        mult_16_res_sva_1 <= z_out_40;
        mult_17_res_sva_1 <= z_out_42;
        mult_18_res_sva_1 <= z_out_44;
        mult_19_res_sva_1 <= z_out_46;
        mult_20_res_sva_1 <= z_out_48;
        mult_21_res_sva_1 <= z_out_55;
        mult_22_res_sva_1 <= z_out_82;
        mult_23_res_sva_1 <= z_out_83;
        mult_24_res_sva_1 <= z_out_84;
        mult_25_res_sva_1 <= mult_25_res_sva_2;
        mult_26_res_sva_1 <= mult_26_res_sva_2;
        mult_27_res_sva_1 <= mult_27_res_sva_2;
        mult_28_res_sva_1 <= mult_28_res_sva_2;
        mult_29_res_sva_1 <= mult_29_res_sva_2;
        mult_30_res_sva_1 <= mult_30_res_sva_2;
        mult_31_res_sva_1 <= mult_31_res_sva_2;
        tmp_30_lpi_3_dfm_8 <= tmp_30_lpi_3_dfm_7;
        tmp_28_lpi_3_dfm_8 <= tmp_28_lpi_3_dfm_7;
        tmp_26_lpi_3_dfm_8 <= tmp_26_lpi_3_dfm_7;
        tmp_24_lpi_3_dfm_8 <= tmp_24_lpi_3_dfm_7;
        tmp_22_lpi_3_dfm_8 <= tmp_22_lpi_3_dfm_7;
        tmp_20_lpi_3_dfm_8 <= tmp_20_lpi_3_dfm_7;
        tmp_18_lpi_3_dfm_8 <= tmp_18_lpi_3_dfm_7;
        tmp_16_lpi_3_dfm_8 <= tmp_16_lpi_3_dfm_7;
        tmp_14_lpi_3_dfm_8 <= tmp_14_lpi_3_dfm_7;
        tmp_12_lpi_3_dfm_8 <= tmp_12_lpi_3_dfm_7;
        tmp_10_lpi_3_dfm_8 <= tmp_10_lpi_3_dfm_7;
        tmp_8_lpi_3_dfm_8 <= tmp_8_lpi_3_dfm_7;
        tmp_6_lpi_3_dfm_8 <= tmp_6_lpi_3_dfm_7;
        tmp_4_lpi_3_dfm_8 <= tmp_4_lpi_3_dfm_7;
        tmp_2_lpi_3_dfm_8 <= tmp_2_lpi_3_dfm_7;
        tmp_lpi_3_dfm_8 <= tmp_lpi_3_dfm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        mult_31_slc_32_svs_st_1 <= '0';
        mult_30_slc_32_svs_st_1 <= '0';
        mult_29_slc_32_svs_st_1 <= '0';
        mult_28_slc_32_svs_st_1 <= '0';
        mult_27_slc_32_svs_st_1 <= '0';
        mult_26_slc_32_svs_st_1 <= '0';
        mult_25_slc_32_svs_st_1 <= '0';
        mult_24_slc_32_svs_st_1 <= '0';
        mult_23_slc_32_svs_st_1 <= '0';
        mult_22_slc_32_svs_st_1 <= '0';
        mult_21_slc_32_svs_st_1 <= '0';
        mult_20_slc_32_svs_st_1 <= '0';
        mult_19_slc_32_svs_st_1 <= '0';
        mult_18_slc_32_svs_st_1 <= '0';
        mult_17_slc_32_svs_st_1 <= '0';
        mult_16_slc_32_svs_st_1 <= '0';
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_9 <= '0';
      ELSIF ( mult_31_if_and_cse = '1' ) THEN
        mult_31_slc_32_svs_st_1 <= mult_31_if_acc_1_nl(32);
        mult_30_slc_32_svs_st_1 <= mult_30_if_acc_1_nl(32);
        mult_29_slc_32_svs_st_1 <= mult_29_if_acc_1_nl(32);
        mult_28_slc_32_svs_st_1 <= mult_28_if_acc_1_nl(32);
        mult_27_slc_32_svs_st_1 <= mult_27_if_acc_1_nl(32);
        mult_26_slc_32_svs_st_1 <= mult_26_if_acc_1_nl(32);
        mult_25_slc_32_svs_st_1 <= mult_25_if_acc_1_nl(32);
        mult_24_slc_32_svs_st_1 <= mult_24_if_acc_1_nl(32);
        mult_23_slc_32_svs_st_1 <= mult_23_if_acc_1_nl(32);
        mult_22_slc_32_svs_st_1 <= mult_22_if_acc_1_nl(32);
        mult_21_slc_32_svs_st_1 <= mult_21_if_acc_1_nl(32);
        mult_20_slc_32_svs_st_1 <= mult_20_if_acc_1_nl(32);
        mult_19_slc_32_svs_st_1 <= mult_19_if_acc_1_nl(32);
        mult_18_slc_32_svs_st_1 <= mult_18_if_acc_1_nl(32);
        mult_17_slc_32_svs_st_1 <= mult_17_if_acc_1_nl(32);
        mult_16_slc_32_svs_st_1 <= mult_16_if_acc_1_nl(32);
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_9 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4302_itm_1 <= '0';
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_1 <= '0';
      ELSIF ( INNER_LOOP2_r_and_3_cse = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4302_itm_1 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4302_itm;
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_1 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND (NOT (fsm_output(4)))) = '1' ) THEN
        operator_33_true_1_lshift_psp_7_4_sva <= z_out_32(7 DOWNTO 4);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4302_itm <= '0';
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm <= '0';
      ELSIF ( INNER_LOOP2_r_and_4_cse = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4302_itm <= INNER_LOOP1_r_INNER_LOOP1_r_and_2_cse(4);
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm <= INNER_LOOP1_r_INNER_LOOP1_r_and_2_cse(0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_31_z_and_cse = '1' ) THEN
        mult_31_z_asn_itm_4 <= mult_31_z_asn_itm_3;
        mult_30_z_asn_itm_4 <= mult_30_z_asn_itm_3;
        mult_29_z_asn_itm_4 <= mult_29_z_asn_itm_3;
        mult_28_z_asn_itm_4 <= mult_28_z_asn_itm_3;
        mult_27_z_asn_itm_4 <= mult_27_z_asn_itm_3;
        mult_26_z_asn_itm_4 <= mult_26_z_asn_itm_3;
        mult_25_z_asn_itm_4 <= mult_25_z_asn_itm_3;
        mult_24_z_asn_itm_4 <= mult_24_z_asn_itm_3;
        mult_23_z_asn_itm_4 <= mult_23_z_asn_itm_3;
        mult_22_z_asn_itm_4 <= mult_22_z_asn_itm_3;
        mult_21_z_asn_itm_4 <= mult_21_z_asn_itm_3;
        mult_20_z_asn_itm_4 <= mult_20_z_asn_itm_3;
        mult_19_z_asn_itm_4 <= mult_19_z_asn_itm_3;
        mult_18_z_asn_itm_4 <= mult_18_z_asn_itm_3;
        mult_17_z_asn_itm_4 <= mult_17_z_asn_itm_3;
        mult_16_z_asn_itm_4 <= mult_16_z_asn_itm_3;
        tmp_30_lpi_3_dfm_7 <= tmp_30_lpi_3_dfm_6;
        tmp_28_lpi_3_dfm_7 <= tmp_28_lpi_3_dfm_6;
        tmp_26_lpi_3_dfm_7 <= tmp_26_lpi_3_dfm_6;
        tmp_24_lpi_3_dfm_7 <= tmp_24_lpi_3_dfm_6;
        tmp_22_lpi_3_dfm_7 <= tmp_22_lpi_3_dfm_6;
        tmp_20_lpi_3_dfm_7 <= tmp_20_lpi_3_dfm_6;
        tmp_18_lpi_3_dfm_7 <= tmp_18_lpi_3_dfm_6;
        tmp_16_lpi_3_dfm_7 <= tmp_16_lpi_3_dfm_6;
        tmp_14_lpi_3_dfm_7 <= tmp_14_lpi_3_dfm_6;
        tmp_12_lpi_3_dfm_7 <= tmp_12_lpi_3_dfm_6;
        tmp_10_lpi_3_dfm_7 <= tmp_10_lpi_3_dfm_6;
        tmp_8_lpi_3_dfm_7 <= tmp_8_lpi_3_dfm_6;
        tmp_6_lpi_3_dfm_7 <= tmp_6_lpi_3_dfm_6;
        tmp_4_lpi_3_dfm_7 <= tmp_4_lpi_3_dfm_6;
        tmp_2_lpi_3_dfm_7 <= tmp_2_lpi_3_dfm_6;
        tmp_lpi_3_dfm_7 <= tmp_lpi_3_dfm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_8 <= '0';
      ELSIF ( mult_31_z_and_cse = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_8 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_10 AND INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_9)
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_10 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_10 AND (NOT INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_9))
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_10 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_9 AND INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_8)
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_9 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_9 AND (NOT INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_8))
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_9 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_31_z_and_1_cse = '1' ) THEN
        mult_31_z_asn_itm_3 <= mult_31_z_asn_itm_2;
        mult_30_z_asn_itm_3 <= mult_30_z_asn_itm_2;
        mult_29_z_asn_itm_3 <= mult_29_z_asn_itm_2;
        mult_28_z_asn_itm_3 <= mult_28_z_asn_itm_2;
        mult_27_z_asn_itm_3 <= mult_27_z_asn_itm_2;
        mult_26_z_asn_itm_3 <= mult_26_z_asn_itm_2;
        mult_25_z_asn_itm_3 <= mult_25_z_asn_itm_2;
        mult_24_z_asn_itm_3 <= mult_24_z_asn_itm_2;
        mult_23_z_asn_itm_3 <= mult_23_z_asn_itm_2;
        mult_22_z_asn_itm_3 <= mult_22_z_asn_itm_2;
        mult_21_z_asn_itm_3 <= mult_21_z_asn_itm_2;
        mult_20_z_asn_itm_3 <= mult_20_z_asn_itm_2;
        mult_19_z_asn_itm_3 <= mult_19_z_asn_itm_2;
        mult_18_z_asn_itm_3 <= mult_18_z_asn_itm_2;
        mult_17_z_asn_itm_3 <= mult_17_z_asn_itm_2;
        mult_16_z_asn_itm_3 <= mult_16_z_asn_itm_2;
        tmp_30_lpi_3_dfm_6 <= tmp_30_lpi_3_dfm_5;
        tmp_28_lpi_3_dfm_6 <= tmp_28_lpi_3_dfm_5;
        tmp_26_lpi_3_dfm_6 <= tmp_26_lpi_3_dfm_5;
        tmp_24_lpi_3_dfm_6 <= tmp_24_lpi_3_dfm_5;
        tmp_22_lpi_3_dfm_6 <= tmp_22_lpi_3_dfm_5;
        tmp_20_lpi_3_dfm_6 <= tmp_20_lpi_3_dfm_5;
        tmp_18_lpi_3_dfm_6 <= tmp_18_lpi_3_dfm_5;
        tmp_16_lpi_3_dfm_6 <= tmp_16_lpi_3_dfm_5;
        tmp_14_lpi_3_dfm_6 <= tmp_14_lpi_3_dfm_5;
        tmp_12_lpi_3_dfm_6 <= tmp_12_lpi_3_dfm_5;
        tmp_10_lpi_3_dfm_6 <= tmp_10_lpi_3_dfm_5;
        tmp_8_lpi_3_dfm_6 <= tmp_8_lpi_3_dfm_5;
        tmp_6_lpi_3_dfm_6 <= tmp_6_lpi_3_dfm_5;
        tmp_4_lpi_3_dfm_6 <= tmp_4_lpi_3_dfm_5;
        tmp_2_lpi_3_dfm_6 <= tmp_2_lpi_3_dfm_5;
        tmp_lpi_3_dfm_6 <= tmp_lpi_3_dfm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_7 <= '0';
      ELSIF ( mult_31_z_and_1_cse = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_7 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_8 AND INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_7)
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_8 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_8 AND (NOT INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_7))
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_8 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_31_z_and_2_cse = '1' ) THEN
        mult_31_z_asn_itm_2 <= mult_15_z_asn_itm_1;
        mult_30_z_asn_itm_2 <= mult_14_z_asn_itm_1;
        mult_29_z_asn_itm_2 <= mult_13_z_asn_itm_1;
        mult_28_z_asn_itm_2 <= mult_12_z_asn_itm_1;
        mult_27_z_asn_itm_2 <= mult_11_z_asn_itm_1;
        mult_26_z_asn_itm_2 <= mult_10_z_asn_itm_1;
        mult_25_z_asn_itm_2 <= mult_9_z_asn_itm_1;
        mult_24_z_asn_itm_2 <= mult_8_z_asn_itm_1;
        mult_23_z_asn_itm_2 <= mult_7_z_asn_itm_1;
        mult_22_z_asn_itm_2 <= mult_6_z_asn_itm_1;
        mult_21_z_asn_itm_2 <= mult_5_z_asn_itm_1;
        mult_20_z_asn_itm_2 <= mult_4_z_asn_itm_1;
        mult_19_z_asn_itm_2 <= mult_3_z_asn_itm_1;
        mult_18_z_asn_itm_2 <= mult_2_z_asn_itm_1;
        mult_17_z_asn_itm_2 <= mult_1_z_asn_itm_1;
        mult_16_z_asn_itm_2 <= mult_z_asn_itm_1;
        tmp_30_lpi_3_dfm_5 <= tmp_30_lpi_3_dfm_4;
        tmp_28_lpi_3_dfm_5 <= tmp_28_lpi_3_dfm_4;
        tmp_26_lpi_3_dfm_5 <= tmp_26_lpi_3_dfm_4;
        tmp_24_lpi_3_dfm_5 <= tmp_24_lpi_3_dfm_4;
        tmp_22_lpi_3_dfm_5 <= tmp_22_lpi_3_dfm_4;
        tmp_20_lpi_3_dfm_5 <= tmp_20_lpi_3_dfm_4;
        tmp_18_lpi_3_dfm_5 <= tmp_18_lpi_3_dfm_4;
        tmp_16_lpi_3_dfm_5 <= tmp_16_lpi_3_dfm_4;
        tmp_14_lpi_3_dfm_5 <= tmp_14_lpi_3_dfm_4;
        tmp_12_lpi_3_dfm_5 <= tmp_12_lpi_3_dfm_4;
        tmp_10_lpi_3_dfm_5 <= tmp_10_lpi_3_dfm_4;
        tmp_8_lpi_3_dfm_5 <= tmp_8_lpi_3_dfm_4;
        tmp_6_lpi_3_dfm_5 <= tmp_6_lpi_3_dfm_4;
        tmp_4_lpi_3_dfm_5 <= tmp_4_lpi_3_dfm_4;
        tmp_2_lpi_3_dfm_5 <= tmp_2_lpi_3_dfm_4;
        tmp_lpi_3_dfm_5 <= tmp_lpi_3_dfm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_6 <= '0';
      ELSIF ( mult_31_z_and_2_cse = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_6 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_7 AND INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_6)
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_7 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_7 AND (NOT INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_6))
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_7 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_6 AND INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_5)
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_6 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_6 AND (NOT INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_5))
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_6 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly1_31_f1_and_4_cse = '1' ) THEN
        tmp_30_lpi_3_dfm_4 <= tmp_30_lpi_3_dfm_3;
        tmp_28_lpi_3_dfm_4 <= tmp_28_lpi_3_dfm_3;
        tmp_26_lpi_3_dfm_4 <= tmp_26_lpi_3_dfm_3;
        tmp_24_lpi_3_dfm_4 <= tmp_24_lpi_3_dfm_3;
        tmp_22_lpi_3_dfm_4 <= tmp_22_lpi_3_dfm_3;
        tmp_20_lpi_3_dfm_4 <= tmp_20_lpi_3_dfm_3;
        tmp_18_lpi_3_dfm_4 <= tmp_18_lpi_3_dfm_3;
        tmp_16_lpi_3_dfm_4 <= tmp_16_lpi_3_dfm_3;
        tmp_14_lpi_3_dfm_4 <= tmp_14_lpi_3_dfm_3;
        tmp_12_lpi_3_dfm_4 <= tmp_12_lpi_3_dfm_3;
        tmp_10_lpi_3_dfm_4 <= tmp_10_lpi_3_dfm_3;
        tmp_8_lpi_3_dfm_4 <= tmp_8_lpi_3_dfm_3;
        tmp_6_lpi_3_dfm_4 <= tmp_6_lpi_3_dfm_3;
        tmp_4_lpi_3_dfm_4 <= tmp_4_lpi_3_dfm_3;
        tmp_2_lpi_3_dfm_4 <= tmp_2_lpi_3_dfm_3;
        tmp_lpi_3_dfm_4 <= tmp_lpi_3_dfm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_5 <= '0';
      ELSIF ( butterFly1_31_f1_and_4_cse = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_5 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_5 AND INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_4)
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_5 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_5 AND (NOT INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_4))
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_5 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly1_31_f1_and_5_cse = '1' ) THEN
        tmp_30_lpi_3_dfm_3 <= tmp_30_lpi_3_dfm_2;
        tmp_28_lpi_3_dfm_3 <= tmp_28_lpi_3_dfm_2;
        tmp_26_lpi_3_dfm_3 <= tmp_26_lpi_3_dfm_2;
        tmp_24_lpi_3_dfm_3 <= tmp_24_lpi_3_dfm_2;
        tmp_22_lpi_3_dfm_3 <= tmp_22_lpi_3_dfm_2;
        tmp_20_lpi_3_dfm_3 <= tmp_20_lpi_3_dfm_2;
        tmp_18_lpi_3_dfm_3 <= tmp_18_lpi_3_dfm_2;
        tmp_16_lpi_3_dfm_3 <= tmp_16_lpi_3_dfm_2;
        tmp_14_lpi_3_dfm_3 <= tmp_14_lpi_3_dfm_2;
        tmp_12_lpi_3_dfm_3 <= tmp_12_lpi_3_dfm_2;
        tmp_10_lpi_3_dfm_3 <= tmp_10_lpi_3_dfm_2;
        tmp_8_lpi_3_dfm_3 <= tmp_8_lpi_3_dfm_2;
        tmp_6_lpi_3_dfm_3 <= tmp_6_lpi_3_dfm_2;
        tmp_4_lpi_3_dfm_3 <= tmp_4_lpi_3_dfm_2;
        tmp_2_lpi_3_dfm_3 <= tmp_2_lpi_3_dfm_2;
        tmp_lpi_3_dfm_3 <= tmp_lpi_3_dfm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_4 <= '0';
      ELSIF ( butterFly1_31_f1_and_5_cse = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_4 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_4 AND INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_3)
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_4 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_4 AND (NOT INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_3))
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_4 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly1_31_f1_and_6_cse = '1' ) THEN
        tmp_30_lpi_3_dfm_2 <= tmp_30_lpi_3_dfm_1;
        tmp_28_lpi_3_dfm_2 <= tmp_28_lpi_3_dfm_1;
        tmp_26_lpi_3_dfm_2 <= tmp_26_lpi_3_dfm_1;
        tmp_24_lpi_3_dfm_2 <= tmp_24_lpi_3_dfm_1;
        tmp_22_lpi_3_dfm_2 <= tmp_22_lpi_3_dfm_1;
        tmp_20_lpi_3_dfm_2 <= tmp_20_lpi_3_dfm_1;
        tmp_18_lpi_3_dfm_2 <= tmp_18_lpi_3_dfm_1;
        tmp_16_lpi_3_dfm_2 <= tmp_16_lpi_3_dfm_1;
        tmp_14_lpi_3_dfm_2 <= tmp_14_lpi_3_dfm_1;
        tmp_12_lpi_3_dfm_2 <= tmp_12_lpi_3_dfm_1;
        tmp_10_lpi_3_dfm_2 <= tmp_10_lpi_3_dfm_1;
        tmp_8_lpi_3_dfm_2 <= tmp_8_lpi_3_dfm_1;
        tmp_6_lpi_3_dfm_2 <= tmp_6_lpi_3_dfm_1;
        tmp_4_lpi_3_dfm_2 <= tmp_4_lpi_3_dfm_1;
        tmp_2_lpi_3_dfm_2 <= tmp_2_lpi_3_dfm_1;
        tmp_lpi_3_dfm_2 <= tmp_lpi_3_dfm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_3 <= '0';
      ELSIF ( butterFly1_31_f1_and_6_cse = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_3 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_3 AND INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_2)
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_3 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_3 AND (NOT INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_2))
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_3 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly1_31_f1_and_7_cse = '1' ) THEN
        tmp_30_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_30_i_qa_d, yt_rsc_1_30_i_qa_d,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_28_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_28_i_qa_d, yt_rsc_1_28_i_qa_d,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_26_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_26_i_qa_d, yt_rsc_1_26_i_qa_d,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_24_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_24_i_qa_d, yt_rsc_1_24_i_qa_d,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_22_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_22_i_qa_d, yt_rsc_1_22_i_qa_d,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_20_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_20_i_qa_d, yt_rsc_1_20_i_qa_d,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_18_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_18_i_qa_d, yt_rsc_1_18_i_qa_d,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_16_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_16_i_qa_d, yt_rsc_1_16_i_qa_d,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_14_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_14_i_qa_d, yt_rsc_1_14_i_qa_d,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_12_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_12_i_qa_d, yt_rsc_1_12_i_qa_d,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_10_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_10_i_qa_d, yt_rsc_1_10_i_qa_d,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_8_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_8_i_qa_d, yt_rsc_1_8_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_6_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_6_i_qa_d, yt_rsc_1_6_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_4_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_4_i_qa_d, yt_rsc_1_4_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_2_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_2_i_qa_d, yt_rsc_1_2_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_lpi_3_dfm_1 <= MUX_v_32_2_2(yt_rsc_0_0_i_qa_d, yt_rsc_1_0_i_qa_d, twiddle_h_rsc_0_0_i_s_raddr_core_4);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_2 <= '0';
      ELSIF ( (core_wen AND INNER_LOOP2_stage_0_2) = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_2 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_2 AND INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_1)
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_2 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0_2 AND (NOT INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm_1))
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_2 <= INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0 AND INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm)
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_20_itm_1 <= INNER_LOOP2_r_9_4_sva_4_0(4
            DOWNTO 1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP2_stage_0 AND (NOT INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_161_itm))
          = '1' ) THEN
        INNER_LOOP2_r_slc_INNER_LOOP2_r_9_4_4_0_4210_itm_1 <= INNER_LOOP2_r_9_4_sva_4_0(4
            DOWNTO 1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        c_1_sva_1 <= '0';
      ELSIF ( (core_wen AND c_or_cse) = '1' ) THEN
        c_1_sva_1 <= MUX_s_1_2_2((operator_20_false_acc_cse_sva(0)), butterFly2_21_tw_butterFly2_21_tw_or_nl,
            fsm_output(8));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_191_itm_12 <= '0';
      ELSIF ( (core_wen AND INNER_LOOP3_stage_0_12) = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_191_itm_12 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_11;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( modulo_add_32_qelse_and_cse = '1' ) THEN
        modulo_add_32_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_32_sva_1, z_out_89,
            z_out_32_1);
        modulo_add_33_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_33_sva_1, z_out_90,
            z_out_1_32);
        modulo_add_34_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_34_sva_1, z_out_91,
            z_out_2_32);
        modulo_add_35_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_35_sva_1, z_out_99,
            z_out_3_32);
        modulo_add_36_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_36_sva_1, z_out_100,
            z_out_4_32);
        modulo_add_37_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_37_sva_1, z_out_98,
            z_out_5_32);
        modulo_add_38_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_38_sva_1, z_out_97,
            z_out_6_32);
        modulo_add_39_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_39_sva_1, z_out_101,
            z_out_7_32);
        modulo_add_40_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_40_sva_1, z_out_34,
            z_out_8_32);
        modulo_add_41_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_41_sva_1, z_out_35,
            z_out_9_32);
        modulo_add_42_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_42_sva_1, z_out_36,
            z_out_10_32);
        modulo_add_43_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_43_sva_1, z_out_63,
            z_out_11_32);
        modulo_add_44_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_44_sva_1, z_out_61,
            z_out_12_32);
        modulo_add_45_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_45_sva_1, z_out_59,
            z_out_13_32);
        modulo_add_46_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_46_sva_1, z_out_57,
            z_out_14_32);
        modulo_add_47_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_47_sva_1, z_out_53,
            z_out_15_32);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_11 <= '0';
      ELSIF ( modulo_add_32_qelse_and_cse = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_11 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_10;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_11 AND (NOT INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_10))
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_321_itm_11 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_416_itm_10;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_11 AND INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_10)
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_337_itm_11 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_432_itm_10;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly2_and_cse = '1' ) THEN
        modulo_add_base_47_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_126_lpi_3_dfm_8)
            + UNSIGNED(mult_47_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_46_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_124_lpi_3_dfm_8)
            + UNSIGNED(mult_46_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_45_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_122_lpi_3_dfm_8)
            + UNSIGNED(mult_45_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_44_sva_1 <= z_out_85;
        modulo_add_base_43_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_118_lpi_3_dfm_8)
            + UNSIGNED(mult_43_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_42_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_116_lpi_3_dfm_8)
            + UNSIGNED(mult_42_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_41_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_114_lpi_3_dfm_8)
            + UNSIGNED(mult_41_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_40_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_112_lpi_3_dfm_8)
            + UNSIGNED(mult_40_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_39_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_110_lpi_3_dfm_8)
            + UNSIGNED(mult_39_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_38_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_108_lpi_3_dfm_8)
            + UNSIGNED(mult_38_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_37_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_106_lpi_3_dfm_8)
            + UNSIGNED(mult_37_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_36_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_104_lpi_3_dfm_8)
            + UNSIGNED(mult_36_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_35_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_102_lpi_3_dfm_8)
            + UNSIGNED(mult_35_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_34_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_100_lpi_3_dfm_8)
            + UNSIGNED(mult_34_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_33_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_98_lpi_3_dfm_8)
            + UNSIGNED(mult_33_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_32_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_96_lpi_3_dfm_8)
            + UNSIGNED(mult_32_res_lpi_3_dfm_mx0), 32));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        modulo_sub_base_32_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_33_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_34_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_35_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_36_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_37_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_38_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_39_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_40_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_41_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_42_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_43_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_44_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_45_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_46_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_47_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_10 <= '0';
      ELSIF ( butterFly2_and_cse = '1' ) THEN
        modulo_sub_base_32_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_96_lpi_3_dfm_8)
            - SIGNED(mult_32_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_33_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_98_lpi_3_dfm_8)
            - SIGNED(mult_33_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_34_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_100_lpi_3_dfm_8)
            - SIGNED(mult_34_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_35_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_102_lpi_3_dfm_8)
            - SIGNED(mult_35_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_36_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_104_lpi_3_dfm_8)
            - SIGNED(mult_36_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_37_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_106_lpi_3_dfm_8)
            - SIGNED(mult_37_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_38_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_108_lpi_3_dfm_8)
            - SIGNED(mult_38_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_39_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_110_lpi_3_dfm_8)
            - SIGNED(mult_39_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_40_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_112_lpi_3_dfm_8)
            - SIGNED(mult_40_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_41_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_114_lpi_3_dfm_8)
            - SIGNED(mult_41_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_42_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_116_lpi_3_dfm_8)
            - SIGNED(mult_42_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_43_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_118_lpi_3_dfm_8)
            - SIGNED(mult_43_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_44_sva_1 <= z_out_86;
        modulo_sub_base_45_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_122_lpi_3_dfm_8)
            - SIGNED(mult_45_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_46_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_124_lpi_3_dfm_8)
            - SIGNED(mult_46_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_47_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_126_lpi_3_dfm_8)
            - SIGNED(mult_47_res_lpi_3_dfm_mx0), 32));
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_10 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_10 AND (NOT INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_9))
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_416_itm_10 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_10 AND INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_9)
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_432_itm_10 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_47_if_and_cse = '1' ) THEN
        mult_32_res_sva_1 <= mult_32_res_sva_2;
        mult_33_res_sva_1 <= mult_33_res_sva_2;
        mult_34_res_sva_1 <= mult_34_res_sva_2;
        mult_35_res_sva_1 <= mult_35_res_sva_2;
        mult_36_res_sva_1 <= mult_36_res_sva_2;
        mult_37_res_sva_1 <= mult_37_res_sva_2;
        mult_38_res_sva_1 <= mult_38_res_sva_2;
        mult_39_res_sva_1 <= mult_39_res_sva_2;
        mult_40_res_sva_1 <= mult_40_res_sva_2;
        mult_41_res_sva_1 <= mult_41_res_sva_2;
        mult_42_res_sva_1 <= mult_42_res_sva_2;
        mult_43_res_sva_1 <= mult_43_res_sva_2;
        mult_44_res_sva_1 <= mult_44_res_sva_2;
        mult_45_res_sva_1 <= mult_45_res_sva_2;
        mult_46_res_sva_1 <= mult_46_res_sva_2;
        mult_47_res_sva_1 <= mult_47_res_sva_2;
        tmp_126_lpi_3_dfm_8 <= tmp_126_lpi_3_dfm_7;
        tmp_124_lpi_3_dfm_8 <= tmp_124_lpi_3_dfm_7;
        tmp_122_lpi_3_dfm_8 <= tmp_122_lpi_3_dfm_7;
        tmp_120_lpi_3_dfm_8 <= tmp_120_lpi_3_dfm_7;
        tmp_118_lpi_3_dfm_8 <= tmp_118_lpi_3_dfm_7;
        tmp_116_lpi_3_dfm_8 <= tmp_116_lpi_3_dfm_7;
        tmp_114_lpi_3_dfm_8 <= tmp_114_lpi_3_dfm_7;
        tmp_112_lpi_3_dfm_8 <= tmp_112_lpi_3_dfm_7;
        tmp_110_lpi_3_dfm_8 <= tmp_110_lpi_3_dfm_7;
        tmp_108_lpi_3_dfm_8 <= tmp_108_lpi_3_dfm_7;
        tmp_106_lpi_3_dfm_8 <= tmp_106_lpi_3_dfm_7;
        tmp_104_lpi_3_dfm_8 <= tmp_104_lpi_3_dfm_7;
        tmp_102_lpi_3_dfm_8 <= tmp_102_lpi_3_dfm_7;
        tmp_100_lpi_3_dfm_8 <= tmp_100_lpi_3_dfm_7;
        tmp_98_lpi_3_dfm_8 <= tmp_98_lpi_3_dfm_7;
        tmp_96_lpi_3_dfm_8 <= tmp_96_lpi_3_dfm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        mult_47_slc_32_svs_st_1 <= '0';
        mult_46_slc_32_svs_st_1 <= '0';
        mult_45_slc_32_svs_st_1 <= '0';
        mult_44_slc_32_svs_st_1 <= '0';
        mult_43_slc_32_svs_st_1 <= '0';
        mult_42_slc_32_svs_st_1 <= '0';
        mult_41_slc_32_svs_st_1 <= '0';
        mult_40_slc_32_svs_st_1 <= '0';
        mult_39_slc_32_svs_st_1 <= '0';
        mult_38_slc_32_svs_st_1 <= '0';
        mult_37_slc_32_svs_st_1 <= '0';
        mult_36_slc_32_svs_st_1 <= '0';
        mult_35_slc_32_svs_st_1 <= '0';
        mult_34_slc_32_svs_st_1 <= '0';
        mult_33_slc_32_svs_st_1 <= '0';
        mult_32_slc_32_svs_st_1 <= '0';
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_9 <= '0';
      ELSIF ( mult_47_if_and_cse = '1' ) THEN
        mult_47_slc_32_svs_st_1 <= z_out_16_32;
        mult_46_slc_32_svs_st_1 <= z_out_17_32;
        mult_45_slc_32_svs_st_1 <= z_out_18_32;
        mult_44_slc_32_svs_st_1 <= z_out_25_32;
        mult_43_slc_32_svs_st_1 <= z_out_19_32;
        mult_42_slc_32_svs_st_1 <= z_out_26_32;
        mult_41_slc_32_svs_st_1 <= z_out_20_32;
        mult_40_slc_32_svs_st_1 <= z_out_27_32;
        mult_39_slc_32_svs_st_1 <= z_out_21_32;
        mult_38_slc_32_svs_st_1 <= z_out_28_32;
        mult_37_slc_32_svs_st_1 <= z_out_22_32;
        mult_36_slc_32_svs_st_1 <= z_out_29_32;
        mult_35_slc_32_svs_st_1 <= z_out_23_32;
        mult_34_slc_32_svs_st_1 <= z_out_30_32;
        mult_33_slc_32_svs_st_1 <= z_out_24_32;
        mult_32_slc_32_svs_st_1 <= z_out_31_32;
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_9 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        butterFly2_15_tw_equal_tmp_1 <= '0';
        butterFly2_15_tw_equal_tmp_3_1 <= '0';
        butterFly2_15_tw_equal_tmp_5_1 <= '0';
        butterFly2_15_tw_equal_tmp_6_1 <= '0';
        butterFly2_15_tw_equal_tmp_7_1 <= '0';
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_1 <= '0';
      ELSIF ( butterFly2_15_tw_and_cse = '1' ) THEN
        butterFly2_15_tw_equal_tmp_1 <= NOT(CONV_SL_1_1(operator_33_true_2_lshift_psp_2_0_sva/=STD_LOGIC_VECTOR'("000")));
        butterFly2_15_tw_equal_tmp_3_1 <= CONV_SL_1_1(operator_33_true_2_lshift_psp_2_0_sva=STD_LOGIC_VECTOR'("011"));
        butterFly2_15_tw_equal_tmp_5_1 <= CONV_SL_1_1(operator_33_true_2_lshift_psp_2_0_sva=STD_LOGIC_VECTOR'("101"));
        butterFly2_15_tw_equal_tmp_6_1 <= CONV_SL_1_1(operator_33_true_2_lshift_psp_2_0_sva=STD_LOGIC_VECTOR'("110"));
        butterFly2_15_tw_equal_tmp_7_1 <= CONV_SL_1_1(operator_33_true_2_lshift_psp_2_0_sva=STD_LOGIC_VECTOR'("111"));
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_1 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_33_true_2_lshift_psp_2_0_sva <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( (core_wen AND (NOT (fsm_output(6)))) = '1' ) THEN
        operator_33_true_2_lshift_psp_2_0_sva <= z_out_32(2 DOWNTO 0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_47_z_and_cse = '1' ) THEN
        mult_47_z_asn_itm_4 <= mult_47_z_asn_itm_3;
        mult_46_z_asn_itm_4 <= mult_46_z_asn_itm_3;
        mult_45_z_asn_itm_4 <= mult_45_z_asn_itm_3;
        mult_44_z_asn_itm_4 <= mult_44_z_asn_itm_3;
        mult_43_z_asn_itm_4 <= mult_43_z_asn_itm_3;
        mult_42_z_asn_itm_4 <= mult_42_z_asn_itm_3;
        mult_41_z_asn_itm_4 <= mult_41_z_asn_itm_3;
        mult_40_z_asn_itm_4 <= mult_40_z_asn_itm_3;
        mult_39_z_asn_itm_4 <= mult_39_z_asn_itm_3;
        mult_38_z_asn_itm_4 <= mult_38_z_asn_itm_3;
        mult_37_z_asn_itm_4 <= mult_37_z_asn_itm_3;
        mult_36_z_asn_itm_4 <= mult_36_z_asn_itm_3;
        mult_35_z_asn_itm_4 <= mult_35_z_asn_itm_3;
        mult_34_z_asn_itm_4 <= mult_34_z_asn_itm_3;
        mult_33_z_asn_itm_4 <= mult_33_z_asn_itm_3;
        mult_32_z_asn_itm_4 <= mult_32_z_asn_itm_3;
        tmp_126_lpi_3_dfm_7 <= tmp_126_lpi_3_dfm_6;
        tmp_124_lpi_3_dfm_7 <= tmp_124_lpi_3_dfm_6;
        tmp_122_lpi_3_dfm_7 <= tmp_122_lpi_3_dfm_6;
        tmp_120_lpi_3_dfm_7 <= tmp_120_lpi_3_dfm_6;
        tmp_118_lpi_3_dfm_7 <= tmp_118_lpi_3_dfm_6;
        tmp_116_lpi_3_dfm_7 <= tmp_116_lpi_3_dfm_6;
        tmp_114_lpi_3_dfm_7 <= tmp_114_lpi_3_dfm_6;
        tmp_112_lpi_3_dfm_7 <= tmp_112_lpi_3_dfm_6;
        tmp_110_lpi_3_dfm_7 <= tmp_110_lpi_3_dfm_6;
        tmp_108_lpi_3_dfm_7 <= tmp_108_lpi_3_dfm_6;
        tmp_106_lpi_3_dfm_7 <= tmp_106_lpi_3_dfm_6;
        tmp_104_lpi_3_dfm_7 <= tmp_104_lpi_3_dfm_6;
        tmp_102_lpi_3_dfm_7 <= tmp_102_lpi_3_dfm_6;
        tmp_100_lpi_3_dfm_7 <= tmp_100_lpi_3_dfm_6;
        tmp_98_lpi_3_dfm_7 <= tmp_98_lpi_3_dfm_6;
        tmp_96_lpi_3_dfm_7 <= tmp_96_lpi_3_dfm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_8 <= '0';
      ELSIF ( mult_47_z_and_cse = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_8 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_9 AND INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_8)
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_9 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_9 AND (NOT INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_8))
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_9 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_8 AND INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_7)
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_8 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_8 AND (NOT INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_7))
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_8 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_47_z_and_1_cse = '1' ) THEN
        mult_47_z_asn_itm_3 <= mult_47_z_asn_itm_2;
        mult_46_z_asn_itm_3 <= mult_46_z_asn_itm_2;
        mult_45_z_asn_itm_3 <= mult_45_z_asn_itm_2;
        mult_44_z_asn_itm_3 <= mult_44_z_asn_itm_2;
        mult_43_z_asn_itm_3 <= mult_43_z_asn_itm_2;
        mult_42_z_asn_itm_3 <= mult_42_z_asn_itm_2;
        mult_41_z_asn_itm_3 <= mult_41_z_asn_itm_2;
        mult_40_z_asn_itm_3 <= mult_40_z_asn_itm_2;
        mult_39_z_asn_itm_3 <= mult_39_z_asn_itm_2;
        mult_38_z_asn_itm_3 <= mult_38_z_asn_itm_2;
        mult_37_z_asn_itm_3 <= mult_37_z_asn_itm_2;
        mult_36_z_asn_itm_3 <= mult_36_z_asn_itm_2;
        mult_35_z_asn_itm_3 <= mult_35_z_asn_itm_2;
        mult_34_z_asn_itm_3 <= mult_34_z_asn_itm_2;
        mult_33_z_asn_itm_3 <= mult_33_z_asn_itm_2;
        mult_32_z_asn_itm_3 <= mult_32_z_asn_itm_2;
        tmp_126_lpi_3_dfm_6 <= tmp_126_lpi_3_dfm_5;
        tmp_124_lpi_3_dfm_6 <= tmp_124_lpi_3_dfm_5;
        tmp_122_lpi_3_dfm_6 <= tmp_122_lpi_3_dfm_5;
        tmp_120_lpi_3_dfm_6 <= tmp_120_lpi_3_dfm_5;
        tmp_118_lpi_3_dfm_6 <= tmp_118_lpi_3_dfm_5;
        tmp_116_lpi_3_dfm_6 <= tmp_116_lpi_3_dfm_5;
        tmp_114_lpi_3_dfm_6 <= tmp_114_lpi_3_dfm_5;
        tmp_112_lpi_3_dfm_6 <= tmp_112_lpi_3_dfm_5;
        tmp_110_lpi_3_dfm_6 <= tmp_110_lpi_3_dfm_5;
        tmp_108_lpi_3_dfm_6 <= tmp_108_lpi_3_dfm_5;
        tmp_106_lpi_3_dfm_6 <= tmp_106_lpi_3_dfm_5;
        tmp_104_lpi_3_dfm_6 <= tmp_104_lpi_3_dfm_5;
        tmp_102_lpi_3_dfm_6 <= tmp_102_lpi_3_dfm_5;
        tmp_100_lpi_3_dfm_6 <= tmp_100_lpi_3_dfm_5;
        tmp_98_lpi_3_dfm_6 <= tmp_98_lpi_3_dfm_5;
        tmp_96_lpi_3_dfm_6 <= tmp_96_lpi_3_dfm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_7 <= '0';
      ELSIF ( mult_47_z_and_1_cse = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_7 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_7 AND INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_6)
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_7 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_7 AND (NOT INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_6))
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_7 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_47_z_and_2_cse = '1' ) THEN
        mult_47_z_asn_itm_2 <= mult_z_asn_itm_1;
        mult_46_z_asn_itm_2 <= mult_14_z_asn_itm_1;
        mult_45_z_asn_itm_2 <= mult_9_z_asn_itm_1;
        mult_44_z_asn_itm_2 <= mult_6_z_asn_itm_1;
        mult_43_z_asn_itm_2 <= mult_1_z_asn_itm_1;
        mult_42_z_asn_itm_2 <= mult_3_z_asn_itm_1;
        mult_41_z_asn_itm_2 <= mult_7_z_asn_itm_1;
        mult_40_z_asn_itm_2 <= mult_11_z_asn_itm_1;
        mult_39_z_asn_itm_2 <= mult_13_z_asn_itm_1;
        mult_38_z_asn_itm_2 <= mult_8_z_asn_itm_1;
        mult_37_z_asn_itm_2 <= mult_5_z_asn_itm_1;
        mult_36_z_asn_itm_2 <= mult_2_z_asn_itm_1;
        mult_35_z_asn_itm_2 <= mult_4_z_asn_itm_1;
        mult_34_z_asn_itm_2 <= mult_10_z_asn_itm_1;
        mult_33_z_asn_itm_2 <= mult_12_z_asn_itm_1;
        mult_32_z_asn_itm_2 <= mult_15_z_asn_itm_1;
        tmp_126_lpi_3_dfm_5 <= tmp_126_lpi_3_dfm_4;
        tmp_124_lpi_3_dfm_5 <= tmp_124_lpi_3_dfm_4;
        tmp_122_lpi_3_dfm_5 <= tmp_122_lpi_3_dfm_4;
        tmp_120_lpi_3_dfm_5 <= tmp_120_lpi_3_dfm_4;
        tmp_118_lpi_3_dfm_5 <= tmp_118_lpi_3_dfm_4;
        tmp_116_lpi_3_dfm_5 <= tmp_116_lpi_3_dfm_4;
        tmp_114_lpi_3_dfm_5 <= tmp_114_lpi_3_dfm_4;
        tmp_112_lpi_3_dfm_5 <= tmp_112_lpi_3_dfm_4;
        tmp_110_lpi_3_dfm_5 <= tmp_110_lpi_3_dfm_4;
        tmp_108_lpi_3_dfm_5 <= tmp_108_lpi_3_dfm_4;
        tmp_106_lpi_3_dfm_5 <= tmp_106_lpi_3_dfm_4;
        tmp_104_lpi_3_dfm_5 <= tmp_104_lpi_3_dfm_4;
        tmp_102_lpi_3_dfm_5 <= tmp_102_lpi_3_dfm_4;
        tmp_100_lpi_3_dfm_5 <= tmp_100_lpi_3_dfm_4;
        tmp_98_lpi_3_dfm_5 <= tmp_98_lpi_3_dfm_4;
        tmp_96_lpi_3_dfm_5 <= tmp_96_lpi_3_dfm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_6 <= '0';
      ELSIF ( mult_47_z_and_2_cse = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_6 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_6 AND INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_5)
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_6 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_6 AND (NOT INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_5))
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_6 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP3_r_and_19_cse = '1' ) THEN
        tmp_126_lpi_3_dfm_4 <= tmp_126_lpi_3_dfm_3;
        tmp_124_lpi_3_dfm_4 <= tmp_124_lpi_3_dfm_3;
        tmp_122_lpi_3_dfm_4 <= tmp_122_lpi_3_dfm_3;
        tmp_120_lpi_3_dfm_4 <= tmp_120_lpi_3_dfm_3;
        tmp_118_lpi_3_dfm_4 <= tmp_118_lpi_3_dfm_3;
        tmp_116_lpi_3_dfm_4 <= tmp_116_lpi_3_dfm_3;
        tmp_114_lpi_3_dfm_4 <= tmp_114_lpi_3_dfm_3;
        tmp_112_lpi_3_dfm_4 <= tmp_112_lpi_3_dfm_3;
        tmp_110_lpi_3_dfm_4 <= tmp_110_lpi_3_dfm_3;
        tmp_108_lpi_3_dfm_4 <= tmp_108_lpi_3_dfm_3;
        tmp_106_lpi_3_dfm_4 <= tmp_106_lpi_3_dfm_3;
        tmp_104_lpi_3_dfm_4 <= tmp_104_lpi_3_dfm_3;
        tmp_102_lpi_3_dfm_4 <= tmp_102_lpi_3_dfm_3;
        tmp_100_lpi_3_dfm_4 <= tmp_100_lpi_3_dfm_3;
        tmp_98_lpi_3_dfm_4 <= tmp_98_lpi_3_dfm_3;
        tmp_96_lpi_3_dfm_4 <= tmp_96_lpi_3_dfm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_5 <= '0';
      ELSIF ( INNER_LOOP3_r_and_19_cse = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_5 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_5 AND INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_4)
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_5 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_5 AND (NOT INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_4))
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_5 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP3_r_and_22_cse = '1' ) THEN
        tmp_126_lpi_3_dfm_3 <= tmp_126_lpi_3_dfm_2;
        tmp_124_lpi_3_dfm_3 <= tmp_124_lpi_3_dfm_2;
        tmp_122_lpi_3_dfm_3 <= tmp_122_lpi_3_dfm_2;
        tmp_120_lpi_3_dfm_3 <= tmp_120_lpi_3_dfm_2;
        tmp_118_lpi_3_dfm_3 <= tmp_118_lpi_3_dfm_2;
        tmp_116_lpi_3_dfm_3 <= tmp_116_lpi_3_dfm_2;
        tmp_114_lpi_3_dfm_3 <= tmp_114_lpi_3_dfm_2;
        tmp_112_lpi_3_dfm_3 <= tmp_112_lpi_3_dfm_2;
        tmp_110_lpi_3_dfm_3 <= tmp_110_lpi_3_dfm_2;
        tmp_108_lpi_3_dfm_3 <= tmp_108_lpi_3_dfm_2;
        tmp_106_lpi_3_dfm_3 <= tmp_106_lpi_3_dfm_2;
        tmp_104_lpi_3_dfm_3 <= tmp_104_lpi_3_dfm_2;
        tmp_102_lpi_3_dfm_3 <= tmp_102_lpi_3_dfm_2;
        tmp_100_lpi_3_dfm_3 <= tmp_100_lpi_3_dfm_2;
        tmp_98_lpi_3_dfm_3 <= tmp_98_lpi_3_dfm_2;
        tmp_96_lpi_3_dfm_3 <= tmp_96_lpi_3_dfm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_4 <= '0';
      ELSIF ( INNER_LOOP3_r_and_22_cse = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_4 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_4 AND INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_3)
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_4 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_4 AND (NOT INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_3))
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_4 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP3_r_and_25_cse = '1' ) THEN
        tmp_126_lpi_3_dfm_2 <= tmp_126_lpi_3_dfm_1;
        tmp_124_lpi_3_dfm_2 <= tmp_124_lpi_3_dfm_1;
        tmp_122_lpi_3_dfm_2 <= tmp_122_lpi_3_dfm_1;
        tmp_120_lpi_3_dfm_2 <= tmp_120_lpi_3_dfm_1;
        tmp_118_lpi_3_dfm_2 <= tmp_118_lpi_3_dfm_1;
        tmp_116_lpi_3_dfm_2 <= tmp_116_lpi_3_dfm_1;
        tmp_114_lpi_3_dfm_2 <= tmp_114_lpi_3_dfm_1;
        tmp_112_lpi_3_dfm_2 <= tmp_112_lpi_3_dfm_1;
        tmp_110_lpi_3_dfm_2 <= tmp_110_lpi_3_dfm_1;
        tmp_108_lpi_3_dfm_2 <= tmp_108_lpi_3_dfm_1;
        tmp_106_lpi_3_dfm_2 <= tmp_106_lpi_3_dfm_1;
        tmp_104_lpi_3_dfm_2 <= tmp_104_lpi_3_dfm_1;
        tmp_102_lpi_3_dfm_2 <= tmp_102_lpi_3_dfm_1;
        tmp_100_lpi_3_dfm_2 <= tmp_100_lpi_3_dfm_1;
        tmp_98_lpi_3_dfm_2 <= tmp_98_lpi_3_dfm_1;
        tmp_96_lpi_3_dfm_2 <= tmp_96_lpi_3_dfm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_3 <= '0';
      ELSIF ( INNER_LOOP3_r_and_25_cse = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_3 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_3 AND INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_2)
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_3 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_3 AND (NOT INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_2))
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_3 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( INNER_LOOP3_r_and_28_cse = '1' ) THEN
        tmp_126_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_30_i_qa_d_mxwt, xt_rsc_1_30_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_124_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_28_i_qa_d_mxwt, xt_rsc_1_28_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_122_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_26_i_qa_d_mxwt, xt_rsc_1_26_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_120_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_24_i_qa_d_mxwt, xt_rsc_1_24_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_118_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_22_i_qa_d_mxwt, xt_rsc_1_22_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_116_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_20_i_qa_d_mxwt, xt_rsc_1_20_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_114_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_18_i_qa_d_mxwt, xt_rsc_1_18_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_112_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_16_i_qa_d_mxwt, xt_rsc_1_16_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_110_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_14_i_qa_d_mxwt, xt_rsc_1_14_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_108_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_12_i_qa_d_mxwt, xt_rsc_1_12_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_106_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_10_i_qa_d_mxwt, xt_rsc_1_10_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_104_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_8_i_qa_d_mxwt, xt_rsc_1_8_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_102_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_6_i_qa_d_mxwt, xt_rsc_1_6_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_100_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_4_i_qa_d_mxwt, xt_rsc_1_4_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_98_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_2_i_qa_d_mxwt, xt_rsc_1_2_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
        tmp_96_lpi_3_dfm_1 <= MUX_v_32_2_2(xt_rsc_0_0_i_qa_d_mxwt, xt_rsc_1_0_i_qa_d_mxwt,
            twiddle_h_rsc_0_0_i_s_raddr_core_4);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_2 <= '0';
      ELSIF ( INNER_LOOP3_r_and_28_cse = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_2 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_2 AND INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_1)
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_2 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0_2 AND (NOT INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm_1))
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_2 <= INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0 AND INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm)
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_20_itm_1 <= INNER_LOOP3_r_9_4_sva_4_0(4
            DOWNTO 1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP3_stage_0 AND (NOT INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm))
          = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_4241_itm_1 <= INNER_LOOP3_r_9_4_sva_4_0(4
            DOWNTO 1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm <= '0';
      ELSIF ( (core_wen AND ((fsm_output(5)) OR (INNER_LOOP3_stage_0 AND (NOT (z_out_33(5)))
          AND (fsm_output(6))))) = '1' ) THEN
        INNER_LOOP3_r_slc_INNER_LOOP3_r_9_4_4_0_192_itm <= (z_out_33(0)) AND (fsm_output(6));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( modulo_add_48_qelse_and_cse = '1' ) THEN
        modulo_add_48_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_48_sva_1, z_out_90,
            z_out_15_32);
        modulo_sub_48_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_48_sva_1(30
            DOWNTO 0))), z_out_79, modulo_sub_base_48_sva_1(31));
        modulo_add_49_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_49_sva_1, z_out_101,
            z_out_14_32);
        modulo_sub_49_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_49_sva_1(30
            DOWNTO 0))), z_out_81, modulo_sub_base_49_sva_1(31));
        modulo_add_50_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_50_sva_1, z_out_91,
            z_out_13_32);
        modulo_sub_50_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_50_sva_1(30
            DOWNTO 0))), z_out_77, modulo_sub_base_50_sva_1(31));
        modulo_add_51_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_51_sva_1, z_out_108,
            z_out_12_32);
        modulo_sub_51_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_51_sva_1(30
            DOWNTO 0))), z_out_75, modulo_sub_base_51_sva_1(31));
        modulo_add_52_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_52_sva_1, z_out_89,
            z_out_11_32);
        modulo_sub_52_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_52_sva_1(30
            DOWNTO 0))), z_out_73, modulo_sub_base_52_sva_1(31));
        modulo_add_53_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_53_sva_1, z_out_109,
            z_out_10_32);
        modulo_sub_53_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_53_sva_1(30
            DOWNTO 0))), z_out_71, modulo_sub_base_53_sva_1(31));
        modulo_add_54_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_54_sva_1, z_out_55,
            z_out_9_32);
        modulo_sub_54_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_54_sva_1(30
            DOWNTO 0))), z_out_69, modulo_sub_base_54_sva_1(31));
        modulo_add_55_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_55_sva_1, z_out_83,
            z_out_8_32);
        modulo_sub_55_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_55_sva_1(30
            DOWNTO 0))), z_out_67, modulo_sub_base_55_sva_1(31));
        modulo_add_56_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_56_sva_1, z_out_84,
            z_out_7_32);
        modulo_sub_56_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_56_sva_1(30
            DOWNTO 0))), z_out_65, modulo_sub_base_56_sva_1(31));
        modulo_add_57_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_57_sva_1, z_out_82,
            z_out_6_32);
        modulo_sub_57_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_57_sva_1(30
            DOWNTO 0))), z_out_49, modulo_sub_base_57_sva_1(31));
        modulo_add_58_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_58_sva_1, z_out_48,
            z_out_5_32);
        modulo_sub_58_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_58_sva_1(30
            DOWNTO 0))), z_out_47, modulo_sub_base_58_sva_1(31));
        modulo_add_59_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_59_sva_1, z_out_46,
            z_out_4_32);
        modulo_sub_59_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_59_sva_1(30
            DOWNTO 0))), z_out_45, modulo_sub_base_59_sva_1(31));
        modulo_add_60_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_60_sva_1, z_out_44,
            z_out_3_32);
        modulo_sub_60_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_60_sva_1(30
            DOWNTO 0))), z_out_43, modulo_sub_base_60_sva_1(31));
        modulo_add_61_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_61_sva_1, z_out_42,
            z_out_2_32);
        modulo_sub_61_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_61_sva_1(30
            DOWNTO 0))), z_out_41, modulo_sub_base_61_sva_1(31));
        modulo_add_62_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_62_sva_1, z_out_40,
            z_out_1_32);
        modulo_sub_62_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_62_sva_1(30
            DOWNTO 0))), z_out_39, modulo_sub_base_62_sva_1(31));
        modulo_add_63_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(modulo_add_base_63_sva_1, z_out_38,
            z_out_32_1);
        modulo_sub_63_qr_lpi_3_dfm_1 <= MUX_v_32_2_2(('0' & (modulo_sub_base_63_sva_1(30
            DOWNTO 0))), z_out_37, modulo_sub_base_63_sva_1(31));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_11 <= '0';
      ELSIF ( modulo_add_48_qelse_and_cse = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_11 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_10;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_11 AND (NOT INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_10))
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_321_itm_11 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_10;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_11 AND INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_10)
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_337_itm_11 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_10;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly2_31_and_cse = '1' ) THEN
        modulo_add_base_63_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_62_lpi_3_dfm_8)
            + UNSIGNED(mult_63_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_62_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_60_lpi_3_dfm_8)
            + UNSIGNED(mult_62_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_61_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_58_lpi_3_dfm_8)
            + UNSIGNED(mult_61_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_60_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_56_lpi_3_dfm_8)
            + UNSIGNED(mult_60_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_59_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_54_lpi_3_dfm_8)
            + UNSIGNED(mult_59_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_58_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_52_lpi_3_dfm_8)
            + UNSIGNED(mult_58_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_57_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_50_lpi_3_dfm_8)
            + UNSIGNED(mult_57_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_56_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_48_lpi_3_dfm_8)
            + UNSIGNED(mult_56_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_55_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_46_lpi_3_dfm_8)
            + UNSIGNED(mult_55_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_54_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_44_lpi_3_dfm_8)
            + UNSIGNED(mult_54_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_53_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_42_lpi_3_dfm_8)
            + UNSIGNED(mult_53_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_52_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_40_lpi_3_dfm_8)
            + UNSIGNED(mult_52_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_51_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_38_lpi_3_dfm_8)
            + UNSIGNED(mult_51_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_50_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_36_lpi_3_dfm_8)
            + UNSIGNED(mult_50_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_49_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_34_lpi_3_dfm_8)
            + UNSIGNED(mult_49_res_lpi_3_dfm_mx0), 32));
        modulo_add_base_48_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(tmp_32_lpi_3_dfm_8)
            + UNSIGNED(mult_48_res_lpi_3_dfm_mx0), 32));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        modulo_sub_base_48_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_49_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_50_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_51_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_52_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_53_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_54_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_55_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_56_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_57_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_58_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_59_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_60_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_61_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_62_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        modulo_sub_base_63_sva_1 <= STD_LOGIC_VECTOR'( "00000000000000000000000000000000");
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_10 <= '0';
      ELSIF ( butterFly2_31_and_cse = '1' ) THEN
        modulo_sub_base_48_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_32_lpi_3_dfm_8)
            - SIGNED(mult_48_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_49_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_34_lpi_3_dfm_8)
            - SIGNED(mult_49_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_50_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_36_lpi_3_dfm_8)
            - SIGNED(mult_50_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_51_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_38_lpi_3_dfm_8)
            - SIGNED(mult_51_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_52_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_40_lpi_3_dfm_8)
            - SIGNED(mult_52_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_53_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_42_lpi_3_dfm_8)
            - SIGNED(mult_53_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_54_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_44_lpi_3_dfm_8)
            - SIGNED(mult_54_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_55_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_46_lpi_3_dfm_8)
            - SIGNED(mult_55_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_56_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_48_lpi_3_dfm_8)
            - SIGNED(mult_56_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_57_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_50_lpi_3_dfm_8)
            - SIGNED(mult_57_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_58_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_52_lpi_3_dfm_8)
            - SIGNED(mult_58_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_59_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_54_lpi_3_dfm_8)
            - SIGNED(mult_59_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_60_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_56_lpi_3_dfm_8)
            - SIGNED(mult_60_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_61_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_58_lpi_3_dfm_8)
            - SIGNED(mult_61_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_62_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_60_lpi_3_dfm_8)
            - SIGNED(mult_62_res_lpi_3_dfm_mx0), 32));
        modulo_sub_base_63_sva_1 <= STD_LOGIC_VECTOR(CONV_SIGNED(SIGNED(tmp_62_lpi_3_dfm_8)
            - SIGNED(mult_63_res_lpi_3_dfm_mx0), 32));
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_10 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_63_if_and_cse = '1' ) THEN
        mult_48_res_sva_1 <= mult_48_res_sva_2;
        mult_49_res_sva_1 <= mult_49_res_sva_2;
        mult_50_res_sva_1 <= mult_50_res_sva_2;
        mult_51_res_sva_1 <= mult_51_res_sva_2;
        mult_52_res_sva_1 <= mult_52_res_sva_2;
        mult_53_res_sva_1 <= mult_53_res_sva_2;
        mult_54_res_sva_1 <= mult_54_res_sva_2;
        mult_55_res_sva_1 <= mult_55_res_sva_2;
        mult_56_res_sva_1 <= mult_56_res_sva_2;
        mult_57_res_sva_1 <= mult_57_res_sva_2;
        mult_58_res_sva_1 <= mult_58_res_sva_2;
        mult_59_res_sva_1 <= mult_59_res_sva_2;
        mult_60_res_sva_1 <= mult_60_res_sva_2;
        mult_61_res_sva_1 <= mult_61_res_sva_2;
        mult_62_res_sva_1 <= mult_62_res_sva_2;
        mult_63_res_sva_1 <= mult_63_res_sva_2;
        tmp_62_lpi_3_dfm_8 <= tmp_62_lpi_3_dfm_7;
        tmp_60_lpi_3_dfm_8 <= tmp_60_lpi_3_dfm_7;
        tmp_58_lpi_3_dfm_8 <= tmp_58_lpi_3_dfm_7;
        tmp_56_lpi_3_dfm_8 <= tmp_56_lpi_3_dfm_7;
        tmp_54_lpi_3_dfm_8 <= tmp_54_lpi_3_dfm_7;
        tmp_52_lpi_3_dfm_8 <= tmp_52_lpi_3_dfm_7;
        tmp_50_lpi_3_dfm_8 <= tmp_50_lpi_3_dfm_7;
        tmp_48_lpi_3_dfm_8 <= tmp_48_lpi_3_dfm_7;
        tmp_46_lpi_3_dfm_8 <= tmp_46_lpi_3_dfm_7;
        tmp_44_lpi_3_dfm_8 <= tmp_44_lpi_3_dfm_7;
        tmp_42_lpi_3_dfm_8 <= tmp_42_lpi_3_dfm_7;
        tmp_40_lpi_3_dfm_8 <= tmp_40_lpi_3_dfm_7;
        tmp_38_lpi_3_dfm_8 <= tmp_38_lpi_3_dfm_7;
        tmp_36_lpi_3_dfm_8 <= tmp_36_lpi_3_dfm_7;
        tmp_34_lpi_3_dfm_8 <= tmp_34_lpi_3_dfm_7;
        tmp_32_lpi_3_dfm_8 <= tmp_32_lpi_3_dfm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        mult_63_slc_32_svs_st_1 <= '0';
        mult_62_slc_32_svs_st_1 <= '0';
        mult_61_slc_32_svs_st_1 <= '0';
        mult_60_slc_32_svs_st_1 <= '0';
        mult_59_slc_32_svs_st_1 <= '0';
        mult_58_slc_32_svs_st_1 <= '0';
        mult_57_slc_32_svs_st_1 <= '0';
        mult_56_slc_32_svs_st_1 <= '0';
        mult_55_slc_32_svs_st_1 <= '0';
        mult_54_slc_32_svs_st_1 <= '0';
        mult_53_slc_32_svs_st_1 <= '0';
        mult_52_slc_32_svs_st_1 <= '0';
        mult_51_slc_32_svs_st_1 <= '0';
        mult_50_slc_32_svs_st_1 <= '0';
        mult_49_slc_32_svs_st_1 <= '0';
        mult_48_slc_32_svs_st_1 <= '0';
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_9 <= '0';
      ELSIF ( mult_63_if_and_cse = '1' ) THEN
        mult_63_slc_32_svs_st_1 <= z_out_31_32;
        mult_62_slc_32_svs_st_1 <= z_out_30_32;
        mult_61_slc_32_svs_st_1 <= z_out_29_32;
        mult_60_slc_32_svs_st_1 <= z_out_28_32;
        mult_59_slc_32_svs_st_1 <= z_out_27_32;
        mult_58_slc_32_svs_st_1 <= z_out_26_32;
        mult_57_slc_32_svs_st_1 <= z_out_25_32;
        mult_56_slc_32_svs_st_1 <= z_out_24_32;
        mult_55_slc_32_svs_st_1 <= z_out_23_32;
        mult_54_slc_32_svs_st_1 <= z_out_22_32;
        mult_53_slc_32_svs_st_1 <= z_out_21_32;
        mult_52_slc_32_svs_st_1 <= z_out_20_32;
        mult_51_slc_32_svs_st_1 <= z_out_19_32;
        mult_50_slc_32_svs_st_1 <= z_out_18_32;
        mult_49_slc_32_svs_st_1 <= z_out_17_32;
        mult_48_slc_32_svs_st_1 <= z_out_16_32;
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_9 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4377_itm_1 <= '0';
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_1 <= '0';
      ELSIF ( INNER_LOOP4_r_and_3_cse = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4377_itm_1 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4377_itm;
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_1 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        operator_33_true_3_lshift_psp_1_0_sva <= STD_LOGIC_VECTOR'( "00");
      ELSIF ( (core_wen AND (NOT (fsm_output(8)))) = '1' ) THEN
        operator_33_true_3_lshift_psp_1_0_sva <= operator_33_true_3_lshift_psp_1_0_sva_mx0w2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4377_itm <= '0';
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm <= '0';
      ELSIF ( INNER_LOOP4_r_and_4_cse = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4377_itm <= INNER_LOOP1_r_INNER_LOOP1_r_and_6_cse(4);
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm <= INNER_LOOP1_r_INNER_LOOP1_r_and_6_cse(0);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_63_z_and_cse = '1' ) THEN
        mult_63_z_asn_itm_4 <= mult_63_z_asn_itm_3;
        mult_62_z_asn_itm_4 <= mult_62_z_asn_itm_3;
        mult_61_z_asn_itm_4 <= mult_61_z_asn_itm_3;
        mult_60_z_asn_itm_4 <= mult_60_z_asn_itm_3;
        mult_59_z_asn_itm_4 <= mult_59_z_asn_itm_3;
        mult_58_z_asn_itm_4 <= mult_58_z_asn_itm_3;
        mult_57_z_asn_itm_4 <= mult_57_z_asn_itm_3;
        mult_56_z_asn_itm_4 <= mult_56_z_asn_itm_3;
        mult_55_z_asn_itm_4 <= mult_55_z_asn_itm_3;
        mult_54_z_asn_itm_4 <= mult_54_z_asn_itm_3;
        mult_53_z_asn_itm_4 <= mult_53_z_asn_itm_3;
        mult_52_z_asn_itm_4 <= mult_52_z_asn_itm_3;
        mult_51_z_asn_itm_4 <= mult_51_z_asn_itm_3;
        mult_50_z_asn_itm_4 <= mult_50_z_asn_itm_3;
        mult_49_z_asn_itm_4 <= mult_49_z_asn_itm_3;
        mult_48_z_asn_itm_4 <= mult_48_z_asn_itm_3;
        tmp_62_lpi_3_dfm_7 <= tmp_62_lpi_3_dfm_6;
        tmp_60_lpi_3_dfm_7 <= tmp_60_lpi_3_dfm_6;
        tmp_58_lpi_3_dfm_7 <= tmp_58_lpi_3_dfm_6;
        tmp_56_lpi_3_dfm_7 <= tmp_56_lpi_3_dfm_6;
        tmp_54_lpi_3_dfm_7 <= tmp_54_lpi_3_dfm_6;
        tmp_52_lpi_3_dfm_7 <= tmp_52_lpi_3_dfm_6;
        tmp_50_lpi_3_dfm_7 <= tmp_50_lpi_3_dfm_6;
        tmp_48_lpi_3_dfm_7 <= tmp_48_lpi_3_dfm_6;
        tmp_46_lpi_3_dfm_7 <= tmp_46_lpi_3_dfm_6;
        tmp_44_lpi_3_dfm_7 <= tmp_44_lpi_3_dfm_6;
        tmp_42_lpi_3_dfm_7 <= tmp_42_lpi_3_dfm_6;
        tmp_40_lpi_3_dfm_7 <= tmp_40_lpi_3_dfm_6;
        tmp_38_lpi_3_dfm_7 <= tmp_38_lpi_3_dfm_6;
        tmp_36_lpi_3_dfm_7 <= tmp_36_lpi_3_dfm_6;
        tmp_34_lpi_3_dfm_7 <= tmp_34_lpi_3_dfm_6;
        tmp_32_lpi_3_dfm_7 <= tmp_32_lpi_3_dfm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_8 <= '0';
      ELSIF ( mult_63_z_and_cse = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_8 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_10 AND INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_9)
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_10 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_10 AND (NOT INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_9))
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_10 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_9;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_9 AND INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_8)
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_9 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_9 AND (NOT INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_8))
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_9 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_8;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_63_z_and_1_cse = '1' ) THEN
        mult_63_z_asn_itm_3 <= mult_63_z_asn_itm_2;
        mult_62_z_asn_itm_3 <= mult_62_z_asn_itm_2;
        mult_61_z_asn_itm_3 <= mult_61_z_asn_itm_2;
        mult_60_z_asn_itm_3 <= mult_60_z_asn_itm_2;
        mult_59_z_asn_itm_3 <= mult_59_z_asn_itm_2;
        mult_58_z_asn_itm_3 <= mult_58_z_asn_itm_2;
        mult_57_z_asn_itm_3 <= mult_57_z_asn_itm_2;
        mult_56_z_asn_itm_3 <= mult_56_z_asn_itm_2;
        mult_55_z_asn_itm_3 <= mult_55_z_asn_itm_2;
        mult_54_z_asn_itm_3 <= mult_54_z_asn_itm_2;
        mult_53_z_asn_itm_3 <= mult_53_z_asn_itm_2;
        mult_52_z_asn_itm_3 <= mult_52_z_asn_itm_2;
        mult_51_z_asn_itm_3 <= mult_51_z_asn_itm_2;
        mult_50_z_asn_itm_3 <= mult_50_z_asn_itm_2;
        mult_49_z_asn_itm_3 <= mult_49_z_asn_itm_2;
        mult_48_z_asn_itm_3 <= mult_48_z_asn_itm_2;
        tmp_62_lpi_3_dfm_6 <= tmp_62_lpi_3_dfm_5;
        tmp_60_lpi_3_dfm_6 <= tmp_60_lpi_3_dfm_5;
        tmp_58_lpi_3_dfm_6 <= tmp_58_lpi_3_dfm_5;
        tmp_56_lpi_3_dfm_6 <= tmp_56_lpi_3_dfm_5;
        tmp_54_lpi_3_dfm_6 <= tmp_54_lpi_3_dfm_5;
        tmp_52_lpi_3_dfm_6 <= tmp_52_lpi_3_dfm_5;
        tmp_50_lpi_3_dfm_6 <= tmp_50_lpi_3_dfm_5;
        tmp_48_lpi_3_dfm_6 <= tmp_48_lpi_3_dfm_5;
        tmp_46_lpi_3_dfm_6 <= tmp_46_lpi_3_dfm_5;
        tmp_44_lpi_3_dfm_6 <= tmp_44_lpi_3_dfm_5;
        tmp_42_lpi_3_dfm_6 <= tmp_42_lpi_3_dfm_5;
        tmp_40_lpi_3_dfm_6 <= tmp_40_lpi_3_dfm_5;
        tmp_38_lpi_3_dfm_6 <= tmp_38_lpi_3_dfm_5;
        tmp_36_lpi_3_dfm_6 <= tmp_36_lpi_3_dfm_5;
        tmp_34_lpi_3_dfm_6 <= tmp_34_lpi_3_dfm_5;
        tmp_32_lpi_3_dfm_6 <= tmp_32_lpi_3_dfm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_7 <= '0';
      ELSIF ( mult_63_z_and_1_cse = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_7 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_8 AND INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_7)
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_8 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_8 AND (NOT INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_7))
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_8 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_7;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( mult_63_z_and_2_cse = '1' ) THEN
        mult_63_z_asn_itm_2 <= mult_13_z_asn_itm_1;
        mult_62_z_asn_itm_2 <= mult_9_z_asn_itm_1;
        mult_61_z_asn_itm_2 <= mult_5_z_asn_itm_1;
        mult_60_z_asn_itm_2 <= mult_1_z_asn_itm_1;
        mult_59_z_asn_itm_2 <= mult_4_z_asn_itm_1;
        mult_58_z_asn_itm_2 <= mult_7_z_asn_itm_1;
        mult_57_z_asn_itm_2 <= mult_12_z_asn_itm_1;
        mult_56_z_asn_itm_2 <= mult_15_z_asn_itm_1;
        mult_55_z_asn_itm_2 <= mult_11_z_asn_itm_1;
        mult_54_z_asn_itm_2 <= mult_3_z_asn_itm_1;
        mult_53_z_asn_itm_2 <= mult_6_z_asn_itm_1;
        mult_52_z_asn_itm_2 <= mult_14_z_asn_itm_1;
        mult_51_z_asn_itm_2 <= mult_10_z_asn_itm_1;
        mult_50_z_asn_itm_2 <= mult_2_z_asn_itm_1;
        mult_49_z_asn_itm_2 <= mult_8_z_asn_itm_1;
        mult_48_z_asn_itm_2 <= mult_z_asn_itm_1;
        tmp_62_lpi_3_dfm_5 <= tmp_62_lpi_3_dfm_4;
        tmp_60_lpi_3_dfm_5 <= tmp_60_lpi_3_dfm_4;
        tmp_58_lpi_3_dfm_5 <= tmp_58_lpi_3_dfm_4;
        tmp_56_lpi_3_dfm_5 <= tmp_56_lpi_3_dfm_4;
        tmp_54_lpi_3_dfm_5 <= tmp_54_lpi_3_dfm_4;
        tmp_52_lpi_3_dfm_5 <= tmp_52_lpi_3_dfm_4;
        tmp_50_lpi_3_dfm_5 <= tmp_50_lpi_3_dfm_4;
        tmp_48_lpi_3_dfm_5 <= tmp_48_lpi_3_dfm_4;
        tmp_46_lpi_3_dfm_5 <= tmp_46_lpi_3_dfm_4;
        tmp_44_lpi_3_dfm_5 <= tmp_44_lpi_3_dfm_4;
        tmp_42_lpi_3_dfm_5 <= tmp_42_lpi_3_dfm_4;
        tmp_40_lpi_3_dfm_5 <= tmp_40_lpi_3_dfm_4;
        tmp_38_lpi_3_dfm_5 <= tmp_38_lpi_3_dfm_4;
        tmp_36_lpi_3_dfm_5 <= tmp_36_lpi_3_dfm_4;
        tmp_34_lpi_3_dfm_5 <= tmp_34_lpi_3_dfm_4;
        tmp_32_lpi_3_dfm_5 <= tmp_32_lpi_3_dfm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_6 <= '0';
      ELSIF ( mult_63_z_and_2_cse = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_6 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_7 AND INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_6)
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_7 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_7 AND (NOT INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_6))
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_7 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_6 AND INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_5)
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_6 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_6 AND (NOT INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_5))
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_6 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_5;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly2_31_f1_and_4_cse = '1' ) THEN
        tmp_62_lpi_3_dfm_4 <= tmp_62_lpi_3_dfm_3;
        tmp_60_lpi_3_dfm_4 <= tmp_60_lpi_3_dfm_3;
        tmp_58_lpi_3_dfm_4 <= tmp_58_lpi_3_dfm_3;
        tmp_56_lpi_3_dfm_4 <= tmp_56_lpi_3_dfm_3;
        tmp_54_lpi_3_dfm_4 <= tmp_54_lpi_3_dfm_3;
        tmp_52_lpi_3_dfm_4 <= tmp_52_lpi_3_dfm_3;
        tmp_50_lpi_3_dfm_4 <= tmp_50_lpi_3_dfm_3;
        tmp_48_lpi_3_dfm_4 <= tmp_48_lpi_3_dfm_3;
        tmp_46_lpi_3_dfm_4 <= tmp_46_lpi_3_dfm_3;
        tmp_44_lpi_3_dfm_4 <= tmp_44_lpi_3_dfm_3;
        tmp_42_lpi_3_dfm_4 <= tmp_42_lpi_3_dfm_3;
        tmp_40_lpi_3_dfm_4 <= tmp_40_lpi_3_dfm_3;
        tmp_38_lpi_3_dfm_4 <= tmp_38_lpi_3_dfm_3;
        tmp_36_lpi_3_dfm_4 <= tmp_36_lpi_3_dfm_3;
        tmp_34_lpi_3_dfm_4 <= tmp_34_lpi_3_dfm_3;
        tmp_32_lpi_3_dfm_4 <= tmp_32_lpi_3_dfm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_5 <= '0';
      ELSIF ( butterFly2_31_f1_and_4_cse = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_5 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_5 AND INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_4)
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_5 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_5 AND (NOT INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_4))
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_5 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_4;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly2_31_f1_and_5_cse = '1' ) THEN
        tmp_62_lpi_3_dfm_3 <= tmp_62_lpi_3_dfm_2;
        tmp_60_lpi_3_dfm_3 <= tmp_60_lpi_3_dfm_2;
        tmp_58_lpi_3_dfm_3 <= tmp_58_lpi_3_dfm_2;
        tmp_56_lpi_3_dfm_3 <= tmp_56_lpi_3_dfm_2;
        tmp_54_lpi_3_dfm_3 <= tmp_54_lpi_3_dfm_2;
        tmp_52_lpi_3_dfm_3 <= tmp_52_lpi_3_dfm_2;
        tmp_50_lpi_3_dfm_3 <= tmp_50_lpi_3_dfm_2;
        tmp_48_lpi_3_dfm_3 <= tmp_48_lpi_3_dfm_2;
        tmp_46_lpi_3_dfm_3 <= tmp_46_lpi_3_dfm_2;
        tmp_44_lpi_3_dfm_3 <= tmp_44_lpi_3_dfm_2;
        tmp_42_lpi_3_dfm_3 <= tmp_42_lpi_3_dfm_2;
        tmp_40_lpi_3_dfm_3 <= tmp_40_lpi_3_dfm_2;
        tmp_38_lpi_3_dfm_3 <= tmp_38_lpi_3_dfm_2;
        tmp_36_lpi_3_dfm_3 <= tmp_36_lpi_3_dfm_2;
        tmp_34_lpi_3_dfm_3 <= tmp_34_lpi_3_dfm_2;
        tmp_32_lpi_3_dfm_3 <= tmp_32_lpi_3_dfm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_4 <= '0';
      ELSIF ( butterFly2_31_f1_and_5_cse = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_4 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_4 AND INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_3)
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_4 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_4 AND (NOT INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_3))
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_4 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( butterFly2_31_f1_and_6_cse = '1' ) THEN
        tmp_62_lpi_3_dfm_2 <= tmp_30_lpi_3_dfm_1;
        tmp_60_lpi_3_dfm_2 <= tmp_28_lpi_3_dfm_1;
        tmp_58_lpi_3_dfm_2 <= tmp_26_lpi_3_dfm_1;
        tmp_56_lpi_3_dfm_2 <= tmp_24_lpi_3_dfm_1;
        tmp_54_lpi_3_dfm_2 <= tmp_22_lpi_3_dfm_1;
        tmp_52_lpi_3_dfm_2 <= tmp_20_lpi_3_dfm_1;
        tmp_50_lpi_3_dfm_2 <= tmp_18_lpi_3_dfm_1;
        tmp_48_lpi_3_dfm_2 <= tmp_16_lpi_3_dfm_1;
        tmp_46_lpi_3_dfm_2 <= tmp_14_lpi_3_dfm_1;
        tmp_44_lpi_3_dfm_2 <= tmp_12_lpi_3_dfm_1;
        tmp_42_lpi_3_dfm_2 <= tmp_10_lpi_3_dfm_1;
        tmp_40_lpi_3_dfm_2 <= tmp_8_lpi_3_dfm_1;
        tmp_38_lpi_3_dfm_2 <= tmp_6_lpi_3_dfm_1;
        tmp_36_lpi_3_dfm_2 <= tmp_4_lpi_3_dfm_1;
        tmp_34_lpi_3_dfm_2 <= tmp_2_lpi_3_dfm_1;
        tmp_32_lpi_3_dfm_2 <= tmp_lpi_3_dfm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_3 <= '0';
      ELSIF ( butterFly2_31_f1_and_6_cse = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_3 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_3 AND INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_2)
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_3 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_3 AND (NOT INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_2))
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_3 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_2 <= '0';
      ELSIF ( (core_wen AND INNER_LOOP4_stage_0_2) = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_2 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_2 AND INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_1)
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_2 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0_2 AND (NOT INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm_1))
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_2 <= INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0 AND INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm)
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_20_itm_1 <= INNER_LOOP4_r_9_4_sva_4_0(4
            DOWNTO 1);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (core_wen AND INNER_LOOP4_stage_0 AND (NOT INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_192_itm))
          = '1' ) THEN
        INNER_LOOP4_r_slc_INNER_LOOP4_r_9_4_4_0_4241_itm_1 <= INNER_LOOP4_r_9_4_sva_4_0(4
            DOWNTO 1);
      END IF;
    END IF;
  END PROCESS;
  INNER_LOOP2_tw_and_nl <= operator_33_true_1_lshift_psp_7_4_sva AND (INNER_LOOP2_r_9_4_sva_4_0(3
      DOWNTO 0));
  nor_4_nl <= NOT((fsm_output(7)) OR (fsm_output(4)) OR (fsm_output(8)));
  modulo_add_20_qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_base_20_sva_1)
      - UNSIGNED(p_sva), 32));
  modulo_add_21_qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_base_21_sva_1)
      - UNSIGNED(p_sva), 32));
  modulo_add_22_qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_base_22_sva_1)
      - UNSIGNED(p_sva), 32));
  modulo_add_23_qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_base_23_sva_1)
      - UNSIGNED(p_sva), 32));
  modulo_add_24_qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_base_24_sva_1)
      - UNSIGNED(p_sva), 32));
  modulo_add_25_qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_base_25_sva_1)
      - UNSIGNED(p_sva), 32));
  modulo_add_26_qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_base_26_sva_1)
      - UNSIGNED(p_sva), 32));
  modulo_add_27_qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_base_27_sva_1)
      - UNSIGNED(p_sva), 32));
  modulo_add_28_qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_base_28_sva_1)
      - UNSIGNED(p_sva), 32));
  modulo_add_29_qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_base_29_sva_1)
      - UNSIGNED(p_sva), 32));
  modulo_add_30_qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_base_30_sva_1)
      - UNSIGNED(p_sva), 32));
  modulo_add_31_qif_acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_base_31_sva_1)
      - UNSIGNED(p_sva), 32));
  mult_31_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_31_res_sva_2)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_30_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_30_res_sva_2)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_29_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_29_res_sva_2)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_28_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_28_res_sva_2)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_27_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_27_res_sva_2)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_26_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_26_res_sva_2)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_25_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_25_res_sva_2)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_24_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & z_out_84)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_23_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & z_out_83)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_22_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & z_out_82)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_21_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & z_out_55)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_20_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & z_out_48)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_19_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & z_out_46)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_18_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & z_out_44)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_17_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & z_out_42)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  mult_16_if_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & z_out_40)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT p_sva), 32), 33) + UNSIGNED'( "000000000000000000000000000000001"),
      33));
  butterFly2_21_tw_butterFly2_21_tw_or_nl <= c_1_sva_1 OR INNER_LOOP4_nor_tmp;
  modulo_add_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_sva_1), (NOT modulo_add_base_16_sva_1),
      (NOT modulo_add_base_32_sva_1), (NOT modulo_add_base_63_sva_1), STD_LOGIC_VECTOR'(
      (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_32_1 <= acc_nl(33);
  modulo_add_1_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_1_sva_1), (NOT
      modulo_add_base_17_sva_1), (NOT modulo_add_base_33_sva_1), (NOT modulo_add_base_62_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_1_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_1_32 <= acc_1_nl(33);
  modulo_add_2_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_2_sva_1), (NOT
      modulo_add_base_18_sva_1), (NOT modulo_add_base_34_sva_1), (NOT modulo_add_base_61_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_2_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_2_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_2_32 <= acc_2_nl(33);
  modulo_add_3_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_3_sva_1), (NOT
      modulo_add_base_19_sva_1), (NOT modulo_add_base_35_sva_1), (NOT modulo_add_base_60_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_3_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_3_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_3_32 <= acc_3_nl(33);
  modulo_add_4_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_4_sva_1), (NOT
      modulo_add_base_20_sva_1), (NOT modulo_add_base_36_sva_1), (NOT modulo_add_base_59_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_4_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_4_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_4_32 <= acc_4_nl(33);
  modulo_add_5_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_5_sva_1), (NOT
      modulo_add_base_21_sva_1), (NOT modulo_add_base_37_sva_1), (NOT modulo_add_base_58_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_5_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_5_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_5_32 <= acc_5_nl(33);
  modulo_add_6_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_6_sva_1), (NOT
      modulo_add_base_22_sva_1), (NOT modulo_add_base_38_sva_1), (NOT modulo_add_base_57_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_6_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_6_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_6_32 <= acc_6_nl(33);
  modulo_add_7_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_7_sva_1), (NOT
      modulo_add_base_23_sva_1), (NOT modulo_add_base_39_sva_1), (NOT modulo_add_base_56_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_7_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_7_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_7_32 <= acc_7_nl(33);
  modulo_add_8_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_8_sva_1), (NOT
      modulo_add_base_24_sva_1), (NOT modulo_add_base_40_sva_1), (NOT modulo_add_base_55_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_8_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_8_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_8_32 <= acc_8_nl(33);
  modulo_add_9_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_9_sva_1), (NOT
      modulo_add_base_25_sva_1), (NOT modulo_add_base_41_sva_1), (NOT modulo_add_base_54_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_9_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_9_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_9_32 <= acc_9_nl(33);
  modulo_add_10_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_10_sva_1), (NOT
      modulo_add_base_26_sva_1), (NOT modulo_add_base_42_sva_1), (NOT modulo_add_base_53_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_10_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_10_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_10_32 <= acc_10_nl(33);
  modulo_add_11_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_11_sva_1), (NOT
      modulo_add_base_27_sva_1), (NOT modulo_add_base_43_sva_1), (NOT modulo_add_base_52_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_11_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_11_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_11_32 <= acc_11_nl(33);
  modulo_add_12_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_12_sva_1), (NOT
      modulo_add_base_28_sva_1), (NOT modulo_add_base_44_sva_1), (NOT modulo_add_base_51_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_12_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_12_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_12_32 <= acc_12_nl(33);
  modulo_add_13_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_13_sva_1), (NOT
      modulo_add_base_29_sva_1), (NOT modulo_add_base_45_sva_1), (NOT modulo_add_base_50_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_13_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_13_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_13_32 <= acc_13_nl(33);
  modulo_add_14_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_14_sva_1), (NOT
      modulo_add_base_30_sva_1), (NOT modulo_add_base_46_sva_1), (NOT modulo_add_base_49_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_14_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_14_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_14_32 <= acc_14_nl(33);
  modulo_add_15_mux1h_3_nl <= MUX1HOT_v_32_4_2((NOT modulo_add_base_15_sva_1), (NOT
      modulo_add_base_31_sva_1), (NOT modulo_add_base_47_sva_1), (NOT modulo_add_base_48_sva_1),
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_15_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & p_sva & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(modulo_add_15_mux1h_3_nl
      & '1'), 33), 34), 34));
  z_out_15_32 <= acc_15_nl(33);
  mult_15_if_mux1h_4_nl <= MUX1HOT_v_32_3_2(mult_15_res_sva_2, mult_47_res_sva_2,
      mult_48_res_sva_2, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_16_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_15_if_mux1h_4_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_16_32 <= acc_16_nl(33);
  mult_14_if_mux1h_4_nl <= MUX1HOT_v_32_3_2(mult_14_res_sva_2, mult_46_res_sva_2,
      mult_49_res_sva_2, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_17_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_14_if_mux1h_4_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_17_32 <= acc_17_nl(33);
  mult_13_if_mux1h_4_nl <= MUX1HOT_v_32_3_2(mult_13_res_sva_2, mult_45_res_sva_2,
      mult_50_res_sva_2, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_18_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_13_if_mux1h_4_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_18_32 <= acc_18_nl(33);
  mult_12_if_mux1h_6_nl <= MUX1HOT_v_32_3_2(mult_12_res_sva_2, mult_43_res_sva_2,
      mult_51_res_sva_2, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_19_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_12_if_mux1h_6_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_19_32 <= acc_19_nl(33);
  mult_11_if_mux1h_4_nl <= MUX1HOT_v_32_3_2(mult_11_res_sva_2, mult_41_res_sva_2,
      mult_52_res_sva_2, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_20_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_11_if_mux1h_4_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_20_32 <= acc_20_nl(33);
  mult_10_if_mux1h_4_nl <= MUX1HOT_v_32_3_2(mult_10_res_sva_2, mult_39_res_sva_2,
      mult_53_res_sva_2, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_21_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_10_if_mux1h_4_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_21_32 <= acc_21_nl(33);
  mult_9_if_mux1h_4_nl <= MUX1HOT_v_32_3_2(mult_9_res_sva_2, mult_37_res_sva_2, mult_54_res_sva_2,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_22_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_9_if_mux1h_4_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_22_32 <= acc_22_nl(33);
  mult_8_if_mux1h_4_nl <= MUX1HOT_v_32_3_2(mult_8_res_sva_2, mult_35_res_sva_2, mult_55_res_sva_2,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_23_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_8_if_mux1h_4_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_23_32 <= acc_23_nl(33);
  mult_7_if_mux1h_4_nl <= MUX1HOT_v_32_3_2(mult_7_res_sva_2, mult_33_res_sva_2, mult_56_res_sva_2,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_24_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_7_if_mux1h_4_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_24_32 <= acc_24_nl(33);
  mult_6_if_mux1h_4_nl <= MUX1HOT_v_32_3_2(mult_6_res_sva_2, mult_44_res_sva_2, mult_57_res_sva_2,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_25_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_6_if_mux1h_4_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_25_32 <= acc_25_nl(33);
  mult_5_if_mux1h_6_nl <= MUX1HOT_v_32_3_2(mult_5_res_sva_2, mult_42_res_sva_2, mult_58_res_sva_2,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_26_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_5_if_mux1h_6_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_26_32 <= acc_26_nl(33);
  mult_4_if_mux1h_4_nl <= MUX1HOT_v_32_3_2(mult_4_res_sva_2, mult_40_res_sva_2, mult_59_res_sva_2,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_27_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_4_if_mux1h_4_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_27_32 <= acc_27_nl(33);
  mult_3_if_mux1h_6_nl <= MUX1HOT_v_32_3_2(mult_3_res_sva_2, mult_38_res_sva_2, mult_60_res_sva_2,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_28_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_3_if_mux1h_6_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_28_32 <= acc_28_nl(33);
  mult_2_if_mux1h_6_nl <= MUX1HOT_v_32_3_2(mult_2_res_sva_2, mult_36_res_sva_2, mult_61_res_sva_2,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_29_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_2_if_mux1h_6_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_29_32 <= acc_29_nl(33);
  mult_1_if_mux1h_4_nl <= MUX1HOT_v_32_3_2(mult_1_res_sva_2, mult_34_res_sva_2, mult_62_res_sva_2,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_30_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_1_if_mux1h_4_nl
      & '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34),
      34));
  z_out_30_32 <= acc_30_nl(33);
  mult_if_mux1h_6_nl <= MUX1HOT_v_32_3_2(mult_res_sva_2, mult_32_res_sva_2, mult_63_res_sva_2,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_31_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & mult_if_mux1h_6_nl &
      '1') + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED((NOT p_sva) & '1'), 33), 34), 34));
  z_out_31_32 <= acc_31_nl(33);
  operator_20_false_1_mux_2_nl <= MUX_v_5_2_2(INNER_LOOP2_r_9_4_sva_4_0, INNER_LOOP3_r_9_4_sva_4_0,
      fsm_output(6));
  z_out_33 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(operator_20_false_1_mux_2_nl),
      6) + UNSIGNED'( "000001"), 6));
  modulo_add_40_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_40_sva_1, mult_15_res_sva_1,
      mult_30_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(6)) & (fsm_output(2)) & (fsm_output(4))));
  acc_33_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_40_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_34 <= acc_33_nl(32 DOWNTO 1);
  modulo_add_41_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_41_sva_1, mult_14_res_sva_1,
      mult_25_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(6)) & (fsm_output(2)) & (fsm_output(4))));
  acc_34_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_41_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_35 <= acc_34_nl(32 DOWNTO 1);
  modulo_add_42_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_42_sva_1, mult_13_res_sva_1,
      mult_26_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(6)) & (fsm_output(2)) & (fsm_output(4))));
  acc_35_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_42_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_36 <= acc_35_nl(32 DOWNTO 1);
  modulo_sub_63_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_63_sva_1(30 DOWNTO
      0)), (modulo_sub_base_15_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_37 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_63_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_add_63_qif_mux_2_nl <= MUX_v_32_2_2(modulo_add_base_63_sva_1, mult_10_res_sva_1,
      fsm_output(2));
  acc_37_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_63_qif_mux_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_38 <= acc_37_nl(32 DOWNTO 1);
  modulo_sub_62_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_62_sva_1(30 DOWNTO
      0)), (modulo_sub_base_14_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_39 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_62_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_add_62_qif_mux_2_nl <= MUX_v_32_2_2(modulo_add_base_62_sva_1, mult_16_z_asn_itm_4,
      fsm_output(4));
  modulo_add_62_qif_mux_3_nl <= MUX_v_32_2_2((NOT p_sva), (NOT reg_mult_z_asn_itm_1_cse),
      fsm_output(4));
  acc_39_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_62_qif_mux_2_nl
      & '1') + UNSIGNED(modulo_add_62_qif_mux_3_nl & '1'), 33));
  z_out_40 <= acc_39_nl(32 DOWNTO 1);
  modulo_sub_61_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_61_sva_1(30 DOWNTO
      0)), (modulo_sub_base_13_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_41 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_61_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_add_61_qif_mux_2_nl <= MUX_v_32_2_2(modulo_add_base_61_sva_1, mult_17_z_asn_itm_4,
      fsm_output(4));
  modulo_add_61_qif_mux_3_nl <= MUX_v_32_2_2((NOT p_sva), (NOT reg_mult_1_z_asn_itm_1_cse),
      fsm_output(4));
  acc_41_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_61_qif_mux_2_nl
      & '1') + UNSIGNED(modulo_add_61_qif_mux_3_nl & '1'), 33));
  z_out_42 <= acc_41_nl(32 DOWNTO 1);
  modulo_sub_60_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_60_sva_1(30 DOWNTO
      0)), (modulo_sub_base_12_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_43 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_60_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_add_60_qif_mux_2_nl <= MUX_v_32_2_2(modulo_add_base_60_sva_1, mult_18_z_asn_itm_4,
      fsm_output(4));
  modulo_add_60_qif_mux_3_nl <= MUX_v_32_2_2((NOT p_sva), (NOT reg_mult_2_z_asn_itm_1_cse),
      fsm_output(4));
  acc_43_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_60_qif_mux_2_nl
      & '1') + UNSIGNED(modulo_add_60_qif_mux_3_nl & '1'), 33));
  z_out_44 <= acc_43_nl(32 DOWNTO 1);
  modulo_sub_59_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_59_sva_1(30 DOWNTO
      0)), (modulo_sub_base_11_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_45 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_59_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_add_59_qif_mux_2_nl <= MUX_v_32_2_2(modulo_add_base_59_sva_1, mult_19_z_asn_itm_4,
      fsm_output(4));
  modulo_add_59_qif_mux_3_nl <= MUX_v_32_2_2((NOT p_sva), (NOT reg_mult_3_z_asn_itm_1_cse),
      fsm_output(4));
  acc_45_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_59_qif_mux_2_nl
      & '1') + UNSIGNED(modulo_add_59_qif_mux_3_nl & '1'), 33));
  z_out_46 <= acc_45_nl(32 DOWNTO 1);
  modulo_sub_58_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_58_sva_1(30 DOWNTO
      0)), (modulo_sub_base_10_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_47 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_58_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_add_58_qif_mux_2_nl <= MUX_v_32_2_2(modulo_add_base_58_sva_1, mult_20_z_asn_itm_4,
      fsm_output(4));
  modulo_add_58_qif_mux_3_nl <= MUX_v_32_2_2((NOT p_sva), (NOT reg_mult_4_z_asn_itm_1_cse),
      fsm_output(4));
  acc_47_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_58_qif_mux_2_nl
      & '1') + UNSIGNED(modulo_add_58_qif_mux_3_nl & '1'), 33));
  z_out_48 <= acc_47_nl(32 DOWNTO 1);
  modulo_sub_57_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_57_sva_1(30 DOWNTO
      0)), (modulo_sub_base_9_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_49 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_57_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_16_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_16_sva_1(30 DOWNTO
      0)), (modulo_sub_base_47_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_50 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_16_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  mult_12_if_mux1h_7_nl <= MUX1HOT_v_32_3_2(mult_12_res_sva_1, mult_31_res_sva_1,
      mult_47_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(4)) & (fsm_output(6))));
  acc_50_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_12_if_mux1h_7_nl & '1')
      + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_51 <= acc_50_nl(32 DOWNTO 1);
  modulo_sub_17_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_17_sva_1(30 DOWNTO
      0)), (modulo_sub_base_46_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_52 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_17_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_add_47_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_47_sva_1, mult_6_res_sva_1,
      mult_27_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(6)) & (fsm_output(2)) & (fsm_output(4))));
  acc_52_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_47_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_53 <= acc_52_nl(32 DOWNTO 1);
  modulo_sub_18_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_18_sva_1(30 DOWNTO
      0)), (modulo_sub_base_45_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_54 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_18_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_add_54_qif_mux_2_nl <= MUX_v_32_2_2(modulo_add_base_54_sva_1, mult_21_z_asn_itm_4,
      fsm_output(4));
  modulo_add_54_qif_mux_3_nl <= MUX_v_32_2_2((NOT p_sva), (NOT reg_mult_5_z_asn_itm_1_cse),
      fsm_output(4));
  acc_54_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_54_qif_mux_2_nl
      & '1') + UNSIGNED(modulo_add_54_qif_mux_3_nl & '1'), 33));
  z_out_55 <= acc_54_nl(32 DOWNTO 1);
  modulo_sub_19_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_19_sva_1(30 DOWNTO
      0)), (modulo_sub_base_44_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_56 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_19_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_add_46_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_46_sva_1, mult_7_res_sva_1,
      mult_29_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(6)) & (fsm_output(2)) & (fsm_output(4))));
  acc_56_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_46_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_57 <= acc_56_nl(32 DOWNTO 1);
  modulo_sub_20_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_20_sva_1(30 DOWNTO
      0)), (modulo_sub_base_43_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_58 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_20_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_add_45_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_45_sva_1, mult_8_res_sva_1,
      mult_24_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(6)) & (fsm_output(2)) & (fsm_output(4))));
  acc_58_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_45_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_59 <= acc_58_nl(32 DOWNTO 1);
  modulo_sub_21_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_21_sva_1(30 DOWNTO
      0)), (modulo_sub_base_42_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_60 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_21_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_add_44_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_44_sva_1, mult_9_res_sva_1,
      mult_23_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(6)) & (fsm_output(2)) & (fsm_output(4))));
  acc_60_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_44_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_61 <= acc_60_nl(32 DOWNTO 1);
  modulo_sub_22_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_22_sva_1(30 DOWNTO
      0)), (modulo_sub_base_41_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_62 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_22_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_add_43_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_43_sva_1, mult_11_res_sva_1,
      mult_28_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(6)) & (fsm_output(2)) & (fsm_output(4))));
  acc_62_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_43_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_63 <= acc_62_nl(32 DOWNTO 1);
  modulo_sub_23_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_23_sva_1(30 DOWNTO
      0)), (modulo_sub_base_40_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_64 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_23_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_56_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_56_sva_1(30 DOWNTO
      0)), (modulo_sub_base_8_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_65 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_56_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_24_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_24_sva_1(30 DOWNTO
      0)), (modulo_sub_base_39_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_66 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_24_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_55_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_55_sva_1(30 DOWNTO
      0)), (modulo_sub_base_7_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_67 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_55_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_25_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_25_sva_1(30 DOWNTO
      0)), (modulo_sub_base_38_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_68 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_25_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_54_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_54_sva_1(30 DOWNTO
      0)), (modulo_sub_base_6_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_69 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_54_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_26_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_26_sva_1(30 DOWNTO
      0)), (modulo_sub_base_37_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_70 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_26_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_53_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_53_sva_1(30 DOWNTO
      0)), (modulo_sub_base_5_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_71 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_53_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_27_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_27_sva_1(30 DOWNTO
      0)), (modulo_sub_base_36_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_72 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_27_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_52_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_52_sva_1(30 DOWNTO
      0)), (modulo_sub_base_4_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_73 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_52_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_28_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_28_sva_1(30 DOWNTO
      0)), (modulo_sub_base_35_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_74 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_28_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_51_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_51_sva_1(30 DOWNTO
      0)), (modulo_sub_base_3_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_75 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_51_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_29_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_29_sva_1(30 DOWNTO
      0)), (modulo_sub_base_34_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_76 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_29_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_50_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_50_sva_1(30 DOWNTO
      0)), (modulo_sub_base_2_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_77 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_50_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_30_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_30_sva_1(30 DOWNTO
      0)), (modulo_sub_base_33_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_78 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_30_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_48_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_48_sva_1(30 DOWNTO
      0)), (modulo_sub_base_1_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_79 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_48_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_31_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_31_sva_1(30 DOWNTO
      0)), (modulo_sub_base_32_sva_1(30 DOWNTO 0)), fsm_output(6));
  z_out_80 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_31_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_sub_49_qif_mux_2_nl <= MUX_v_31_2_2((modulo_sub_base_49_sva_1(30 DOWNTO
      0)), (modulo_sub_base_sva_1(30 DOWNTO 0)), fsm_output(2));
  z_out_81 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & modulo_sub_49_qif_mux_2_nl)
      + UNSIGNED(p_sva), 32));
  modulo_add_57_qif_mux_2_nl <= MUX_v_32_2_2(modulo_add_base_57_sva_1, mult_22_z_asn_itm_4,
      fsm_output(4));
  modulo_add_57_qif_mux_3_nl <= MUX_v_32_2_2((NOT p_sva), (NOT reg_mult_6_z_asn_itm_1_cse),
      fsm_output(4));
  acc_81_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_57_qif_mux_2_nl
      & '1') + UNSIGNED(modulo_add_57_qif_mux_3_nl & '1'), 33));
  z_out_82 <= acc_81_nl(32 DOWNTO 1);
  modulo_add_55_qif_mux_2_nl <= MUX_v_32_2_2(modulo_add_base_55_sva_1, mult_23_z_asn_itm_4,
      fsm_output(4));
  modulo_add_55_qif_mux_3_nl <= MUX_v_32_2_2((NOT p_sva), (NOT reg_mult_7_z_asn_itm_1_cse),
      fsm_output(4));
  acc_82_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_55_qif_mux_2_nl
      & '1') + UNSIGNED(modulo_add_55_qif_mux_3_nl & '1'), 33));
  z_out_83 <= acc_82_nl(32 DOWNTO 1);
  modulo_add_56_qif_mux_2_nl <= MUX_v_32_2_2(modulo_add_base_56_sva_1, mult_24_z_asn_itm_4,
      fsm_output(4));
  modulo_add_56_qif_mux_3_nl <= MUX_v_32_2_2((NOT p_sva), (NOT reg_mult_8_z_asn_itm_1_cse),
      fsm_output(4));
  acc_83_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_56_qif_mux_2_nl
      & '1') + UNSIGNED(modulo_add_56_qif_mux_3_nl & '1'), 33));
  z_out_84 <= acc_83_nl(32 DOWNTO 1);
  butterFly1_10_mux_7_cse <= MUX_v_32_2_2(tmp_84_lpi_3_dfm_8, tmp_120_lpi_3_dfm_8,
      fsm_output(6));
  butterFly1_10_mux_8_nl <= MUX_v_32_2_2(mult_10_res_lpi_3_dfm_mx0, mult_44_res_lpi_3_dfm_mx0,
      fsm_output(6));
  z_out_85 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(butterFly1_10_mux_7_cse) +
      UNSIGNED(butterFly1_10_mux_8_nl), 32));
  butterFly1_10_mux_10_nl <= MUX_v_32_2_2((NOT mult_10_res_lpi_3_dfm_mx0), (NOT mult_44_res_lpi_3_dfm_mx0),
      fsm_output(6));
  acc_85_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(butterFly1_10_mux_7_cse &
      '1') + UNSIGNED(butterFly1_10_mux_10_nl & '1'), 33));
  z_out_86 <= acc_85_nl(32 DOWNTO 1);
  modulo_add_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_sva_1, mult_32_res_sva_1,
      mult_48_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_86_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_87 <= acc_86_nl(32 DOWNTO 1);
  modulo_add_1_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_1_sva_1, mult_33_res_sva_1,
      mult_49_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_87_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_1_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_88 <= acc_87_nl(32 DOWNTO 1);
  modulo_add_2_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(modulo_add_base_2_sva_1, modulo_add_base_16_sva_1,
      modulo_add_base_32_sva_1, modulo_add_base_52_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_88_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_2_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_89 <= acc_88_nl(32 DOWNTO 1);
  modulo_add_3_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(modulo_add_base_3_sva_1, modulo_add_base_17_sva_1,
      modulo_add_base_33_sva_1, modulo_add_base_48_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_89_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_3_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_90 <= acc_89_nl(32 DOWNTO 1);
  modulo_add_4_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(modulo_add_base_4_sva_1, modulo_add_base_18_sva_1,
      modulo_add_base_34_sva_1, modulo_add_base_50_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_90_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_4_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_91 <= acc_90_nl(32 DOWNTO 1);
  modulo_add_5_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_5_sva_1, mult_34_res_sva_1,
      mult_50_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_91_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_5_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_92 <= acc_91_nl(32 DOWNTO 1);
  modulo_add_6_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_6_sva_1, mult_35_res_sva_1,
      mult_51_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_92_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_6_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_93 <= acc_92_nl(32 DOWNTO 1);
  modulo_add_7_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_7_sva_1, mult_36_res_sva_1,
      mult_52_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_93_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_7_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_94 <= acc_93_nl(32 DOWNTO 1);
  modulo_add_8_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_8_sva_1, mult_37_res_sva_1,
      mult_53_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_94_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_8_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_95 <= acc_94_nl(32 DOWNTO 1);
  modulo_add_9_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_9_sva_1, mult_38_res_sva_1,
      mult_54_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_95_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_9_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_96 <= acc_95_nl(32 DOWNTO 1);
  modulo_add_10_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_10_sva_1, modulo_add_base_38_sva_1,
      mult_55_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_96_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_10_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_97 <= acc_96_nl(32 DOWNTO 1);
  modulo_add_11_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_11_sva_1, modulo_add_base_37_sva_1,
      mult_56_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_97_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_11_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_98 <= acc_97_nl(32 DOWNTO 1);
  modulo_add_12_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_12_sva_1, modulo_add_base_35_sva_1,
      mult_57_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_98_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_12_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_99 <= acc_98_nl(32 DOWNTO 1);
  modulo_add_13_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_13_sva_1, modulo_add_base_36_sva_1,
      mult_58_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_99_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_13_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_100 <= acc_99_nl(32 DOWNTO 1);
  modulo_add_14_qif_mux1h_2_nl <= MUX1HOT_v_32_4_2(modulo_add_base_14_sva_1, modulo_add_base_19_sva_1,
      modulo_add_base_39_sva_1, modulo_add_base_49_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2))
      & (fsm_output(4)) & (fsm_output(6)) & (fsm_output(8))));
  acc_100_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_14_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_101 <= acc_100_nl(32 DOWNTO 1);
  modulo_add_15_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_15_sva_1, mult_43_res_sva_1,
      mult_59_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_101_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_15_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_102 <= acc_101_nl(32 DOWNTO 1);
  mult_5_if_mux1h_7_nl <= MUX1HOT_v_32_3_2(mult_5_res_sva_1, mult_41_res_sva_1, mult_60_res_sva_1,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_102_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_5_if_mux1h_7_nl & '1')
      + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_103 <= acc_102_nl(32 DOWNTO 1);
  mult_3_if_mux1h_7_nl <= MUX1HOT_v_32_3_2(mult_3_res_sva_1, mult_39_res_sva_1, mult_61_res_sva_1,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_103_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_3_if_mux1h_7_nl & '1')
      + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_104 <= acc_103_nl(32 DOWNTO 1);
  mult_if_mux1h_7_nl <= MUX1HOT_v_32_3_2(mult_res_sva_1, mult_46_res_sva_1, mult_62_res_sva_1,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_104_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_if_mux1h_7_nl & '1')
      + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_105 <= acc_104_nl(32 DOWNTO 1);
  mult_16_if_mux_2_nl <= MUX_v_32_2_2(mult_16_res_sva_1, mult_44_res_sva_1, fsm_output(6));
  acc_105_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_16_if_mux_2_nl & '1')
      + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_106 <= acc_105_nl(32 DOWNTO 1);
  mult_2_if_mux1h_7_nl <= MUX1HOT_v_32_3_2(mult_2_res_sva_1, mult_45_res_sva_1, mult_63_res_sva_1,
      STD_LOGIC_VECTOR'( (fsm_output(2)) & (fsm_output(6)) & (fsm_output(8))));
  acc_106_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(mult_2_if_mux1h_7_nl & '1')
      + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_107 <= acc_106_nl(32 DOWNTO 1);
  modulo_add_51_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_51_sva_1, mult_4_res_sva_1,
      mult_42_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(8)) & (fsm_output(2)) & (fsm_output(6))));
  acc_107_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_51_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_108 <= acc_107_nl(32 DOWNTO 1);
  modulo_add_53_qif_mux1h_2_nl <= MUX1HOT_v_32_3_2(modulo_add_base_53_sva_1, mult_1_res_sva_1,
      mult_40_res_sva_1, STD_LOGIC_VECTOR'( (fsm_output(8)) & (fsm_output(2)) & (fsm_output(6))));
  acc_108_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(modulo_add_53_qif_mux1h_2_nl
      & '1') + UNSIGNED((NOT p_sva) & '1'), 33));
  z_out_109 <= acc_108_nl(32 DOWNTO 1);
END v29;

-- ------------------------------------------------------------------
--  Design Unit:    peaseNTT
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.amba_comps.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;
USE work.ccs_in_pkg_v1.ALL;
USE work.mgc_comps.ALL;
USE work.mgc_shift_comps_v5.ALL;
USE work.BLOCK_2R1W_RBW_pkg.ALL;


ENTITY peaseNTT IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    xt_rsc_0_0_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_0_wea : OUT STD_LOGIC;
    xt_rsc_0_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    xt_rsc_0_1_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_1_wea : OUT STD_LOGIC;
    xt_rsc_0_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    xt_rsc_0_2_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_2_wea : OUT STD_LOGIC;
    xt_rsc_0_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    xt_rsc_0_3_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_3_wea : OUT STD_LOGIC;
    xt_rsc_0_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    xt_rsc_0_4_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_4_wea : OUT STD_LOGIC;
    xt_rsc_0_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    xt_rsc_0_5_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_5_wea : OUT STD_LOGIC;
    xt_rsc_0_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    xt_rsc_0_6_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_6_wea : OUT STD_LOGIC;
    xt_rsc_0_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    xt_rsc_0_7_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_7_wea : OUT STD_LOGIC;
    xt_rsc_0_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    xt_rsc_0_8_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_8_wea : OUT STD_LOGIC;
    xt_rsc_0_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    xt_rsc_0_9_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_9_wea : OUT STD_LOGIC;
    xt_rsc_0_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    xt_rsc_0_10_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_10_wea : OUT STD_LOGIC;
    xt_rsc_0_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    xt_rsc_0_11_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_11_wea : OUT STD_LOGIC;
    xt_rsc_0_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    xt_rsc_0_12_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_12_wea : OUT STD_LOGIC;
    xt_rsc_0_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    xt_rsc_0_13_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_13_wea : OUT STD_LOGIC;
    xt_rsc_0_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    xt_rsc_0_14_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_14_wea : OUT STD_LOGIC;
    xt_rsc_0_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    xt_rsc_0_15_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_15_wea : OUT STD_LOGIC;
    xt_rsc_0_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    xt_rsc_0_16_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_16_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_16_wea : OUT STD_LOGIC;
    xt_rsc_0_16_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_16_lz : OUT STD_LOGIC;
    xt_rsc_0_17_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_17_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_17_wea : OUT STD_LOGIC;
    xt_rsc_0_17_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_17_lz : OUT STD_LOGIC;
    xt_rsc_0_18_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_18_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_18_wea : OUT STD_LOGIC;
    xt_rsc_0_18_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_18_lz : OUT STD_LOGIC;
    xt_rsc_0_19_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_19_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_19_wea : OUT STD_LOGIC;
    xt_rsc_0_19_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_19_lz : OUT STD_LOGIC;
    xt_rsc_0_20_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_20_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_20_wea : OUT STD_LOGIC;
    xt_rsc_0_20_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_20_lz : OUT STD_LOGIC;
    xt_rsc_0_21_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_21_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_21_wea : OUT STD_LOGIC;
    xt_rsc_0_21_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_21_lz : OUT STD_LOGIC;
    xt_rsc_0_22_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_22_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_22_wea : OUT STD_LOGIC;
    xt_rsc_0_22_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_22_lz : OUT STD_LOGIC;
    xt_rsc_0_23_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_23_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_23_wea : OUT STD_LOGIC;
    xt_rsc_0_23_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_23_lz : OUT STD_LOGIC;
    xt_rsc_0_24_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_24_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_24_wea : OUT STD_LOGIC;
    xt_rsc_0_24_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_24_lz : OUT STD_LOGIC;
    xt_rsc_0_25_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_25_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_25_wea : OUT STD_LOGIC;
    xt_rsc_0_25_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_25_lz : OUT STD_LOGIC;
    xt_rsc_0_26_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_26_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_26_wea : OUT STD_LOGIC;
    xt_rsc_0_26_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_26_lz : OUT STD_LOGIC;
    xt_rsc_0_27_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_27_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_27_wea : OUT STD_LOGIC;
    xt_rsc_0_27_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_27_lz : OUT STD_LOGIC;
    xt_rsc_0_28_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_28_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_28_wea : OUT STD_LOGIC;
    xt_rsc_0_28_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_28_lz : OUT STD_LOGIC;
    xt_rsc_0_29_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_29_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_29_wea : OUT STD_LOGIC;
    xt_rsc_0_29_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_29_lz : OUT STD_LOGIC;
    xt_rsc_0_30_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_30_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_30_wea : OUT STD_LOGIC;
    xt_rsc_0_30_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_30_lz : OUT STD_LOGIC;
    xt_rsc_0_31_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_0_31_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_0_31_wea : OUT STD_LOGIC;
    xt_rsc_0_31_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_0_31_lz : OUT STD_LOGIC;
    xt_rsc_1_0_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_0_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_0_wea : OUT STD_LOGIC;
    xt_rsc_1_0_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_0_lz : OUT STD_LOGIC;
    xt_rsc_1_1_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_1_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_1_wea : OUT STD_LOGIC;
    xt_rsc_1_1_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_1_lz : OUT STD_LOGIC;
    xt_rsc_1_2_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_2_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_2_wea : OUT STD_LOGIC;
    xt_rsc_1_2_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_2_lz : OUT STD_LOGIC;
    xt_rsc_1_3_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_3_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_3_wea : OUT STD_LOGIC;
    xt_rsc_1_3_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_3_lz : OUT STD_LOGIC;
    xt_rsc_1_4_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_4_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_4_wea : OUT STD_LOGIC;
    xt_rsc_1_4_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_4_lz : OUT STD_LOGIC;
    xt_rsc_1_5_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_5_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_5_wea : OUT STD_LOGIC;
    xt_rsc_1_5_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_5_lz : OUT STD_LOGIC;
    xt_rsc_1_6_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_6_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_6_wea : OUT STD_LOGIC;
    xt_rsc_1_6_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_6_lz : OUT STD_LOGIC;
    xt_rsc_1_7_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_7_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_7_wea : OUT STD_LOGIC;
    xt_rsc_1_7_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_7_lz : OUT STD_LOGIC;
    xt_rsc_1_8_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_8_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_8_wea : OUT STD_LOGIC;
    xt_rsc_1_8_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_8_lz : OUT STD_LOGIC;
    xt_rsc_1_9_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_9_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_9_wea : OUT STD_LOGIC;
    xt_rsc_1_9_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_9_lz : OUT STD_LOGIC;
    xt_rsc_1_10_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_10_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_10_wea : OUT STD_LOGIC;
    xt_rsc_1_10_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_10_lz : OUT STD_LOGIC;
    xt_rsc_1_11_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_11_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_11_wea : OUT STD_LOGIC;
    xt_rsc_1_11_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_11_lz : OUT STD_LOGIC;
    xt_rsc_1_12_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_12_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_12_wea : OUT STD_LOGIC;
    xt_rsc_1_12_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_12_lz : OUT STD_LOGIC;
    xt_rsc_1_13_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_13_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_13_wea : OUT STD_LOGIC;
    xt_rsc_1_13_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_13_lz : OUT STD_LOGIC;
    xt_rsc_1_14_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_14_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_14_wea : OUT STD_LOGIC;
    xt_rsc_1_14_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_14_lz : OUT STD_LOGIC;
    xt_rsc_1_15_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_15_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_15_wea : OUT STD_LOGIC;
    xt_rsc_1_15_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_15_lz : OUT STD_LOGIC;
    xt_rsc_1_16_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_16_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_16_wea : OUT STD_LOGIC;
    xt_rsc_1_16_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_16_lz : OUT STD_LOGIC;
    xt_rsc_1_17_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_17_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_17_wea : OUT STD_LOGIC;
    xt_rsc_1_17_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_17_lz : OUT STD_LOGIC;
    xt_rsc_1_18_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_18_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_18_wea : OUT STD_LOGIC;
    xt_rsc_1_18_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_18_lz : OUT STD_LOGIC;
    xt_rsc_1_19_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_19_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_19_wea : OUT STD_LOGIC;
    xt_rsc_1_19_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_19_lz : OUT STD_LOGIC;
    xt_rsc_1_20_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_20_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_20_wea : OUT STD_LOGIC;
    xt_rsc_1_20_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_20_lz : OUT STD_LOGIC;
    xt_rsc_1_21_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_21_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_21_wea : OUT STD_LOGIC;
    xt_rsc_1_21_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_21_lz : OUT STD_LOGIC;
    xt_rsc_1_22_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_22_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_22_wea : OUT STD_LOGIC;
    xt_rsc_1_22_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_22_lz : OUT STD_LOGIC;
    xt_rsc_1_23_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_23_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_23_wea : OUT STD_LOGIC;
    xt_rsc_1_23_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_23_lz : OUT STD_LOGIC;
    xt_rsc_1_24_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_24_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_24_wea : OUT STD_LOGIC;
    xt_rsc_1_24_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_24_lz : OUT STD_LOGIC;
    xt_rsc_1_25_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_25_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_25_wea : OUT STD_LOGIC;
    xt_rsc_1_25_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_25_lz : OUT STD_LOGIC;
    xt_rsc_1_26_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_26_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_26_wea : OUT STD_LOGIC;
    xt_rsc_1_26_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_26_lz : OUT STD_LOGIC;
    xt_rsc_1_27_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_27_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_27_wea : OUT STD_LOGIC;
    xt_rsc_1_27_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_27_lz : OUT STD_LOGIC;
    xt_rsc_1_28_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_28_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_28_wea : OUT STD_LOGIC;
    xt_rsc_1_28_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_28_lz : OUT STD_LOGIC;
    xt_rsc_1_29_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_29_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_29_wea : OUT STD_LOGIC;
    xt_rsc_1_29_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_29_lz : OUT STD_LOGIC;
    xt_rsc_1_30_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_30_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_30_wea : OUT STD_LOGIC;
    xt_rsc_1_30_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_30_lz : OUT STD_LOGIC;
    xt_rsc_1_31_adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
    xt_rsc_1_31_da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_1_31_wea : OUT STD_LOGIC;
    xt_rsc_1_31_qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    xt_rsc_triosy_1_31_lz : OUT STD_LOGIC;
    p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    p_rsc_triosy_lz : OUT STD_LOGIC;
    r_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    r_rsc_triosy_lz : OUT STD_LOGIC;
    twiddle_rsc_0_0_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_0_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_0_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_0_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_0_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_0_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_RID : OUT STD_LOGIC;
    twiddle_rsc_0_0_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_0_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_0_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_0_ARID : IN STD_LOGIC;
    twiddle_rsc_0_0_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_0_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_0_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_0_BID : OUT STD_LOGIC;
    twiddle_rsc_0_0_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_0_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_0_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_0_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_0_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_0_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_0_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_0_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_0_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_rsc_0_1_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_1_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_1_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_1_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_1_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_1_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_1_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_1_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_RID : OUT STD_LOGIC;
    twiddle_rsc_0_1_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_1_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_1_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_1_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_1_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_1_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_1_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_1_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_1_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_1_ARID : IN STD_LOGIC;
    twiddle_rsc_0_1_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_1_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_1_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_1_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_1_BID : OUT STD_LOGIC;
    twiddle_rsc_0_1_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_1_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_1_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_1_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_1_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_1_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_1_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_1_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_1_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_1_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_1_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_1_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_1_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_1_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_1_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_1_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_rsc_0_2_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_2_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_2_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_2_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_2_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_2_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_2_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_2_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_RID : OUT STD_LOGIC;
    twiddle_rsc_0_2_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_2_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_2_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_2_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_2_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_2_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_2_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_2_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_2_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_2_ARID : IN STD_LOGIC;
    twiddle_rsc_0_2_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_2_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_2_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_2_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_2_BID : OUT STD_LOGIC;
    twiddle_rsc_0_2_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_2_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_2_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_2_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_2_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_2_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_2_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_2_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_2_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_2_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_2_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_2_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_2_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_2_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_2_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_2_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_rsc_0_3_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_3_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_3_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_3_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_3_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_3_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_3_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_3_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_RID : OUT STD_LOGIC;
    twiddle_rsc_0_3_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_3_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_3_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_3_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_3_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_3_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_3_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_3_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_3_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_3_ARID : IN STD_LOGIC;
    twiddle_rsc_0_3_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_3_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_3_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_3_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_3_BID : OUT STD_LOGIC;
    twiddle_rsc_0_3_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_3_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_3_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_3_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_3_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_3_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_3_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_3_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_3_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_3_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_3_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_3_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_3_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_3_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_3_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_3_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_rsc_0_4_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_4_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_4_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_4_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_4_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_4_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_4_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_4_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_RID : OUT STD_LOGIC;
    twiddle_rsc_0_4_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_4_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_4_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_4_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_4_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_4_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_4_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_4_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_4_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_4_ARID : IN STD_LOGIC;
    twiddle_rsc_0_4_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_4_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_4_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_4_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_4_BID : OUT STD_LOGIC;
    twiddle_rsc_0_4_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_4_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_4_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_4_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_4_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_4_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_4_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_4_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_4_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_4_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_4_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_4_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_4_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_4_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_4_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_4_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_rsc_0_5_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_5_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_5_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_5_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_5_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_5_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_5_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_5_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_RID : OUT STD_LOGIC;
    twiddle_rsc_0_5_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_5_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_5_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_5_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_5_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_5_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_5_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_5_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_5_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_5_ARID : IN STD_LOGIC;
    twiddle_rsc_0_5_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_5_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_5_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_5_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_5_BID : OUT STD_LOGIC;
    twiddle_rsc_0_5_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_5_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_5_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_5_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_5_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_5_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_5_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_5_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_5_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_5_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_5_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_5_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_5_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_5_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_5_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_5_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_rsc_0_6_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_6_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_6_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_6_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_6_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_6_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_6_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_6_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_RID : OUT STD_LOGIC;
    twiddle_rsc_0_6_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_6_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_6_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_6_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_6_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_6_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_6_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_6_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_6_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_6_ARID : IN STD_LOGIC;
    twiddle_rsc_0_6_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_6_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_6_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_6_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_6_BID : OUT STD_LOGIC;
    twiddle_rsc_0_6_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_6_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_6_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_6_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_6_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_6_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_6_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_6_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_6_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_6_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_6_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_6_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_6_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_6_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_6_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_6_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_rsc_0_7_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_7_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_7_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_7_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_7_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_7_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_7_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_7_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_RID : OUT STD_LOGIC;
    twiddle_rsc_0_7_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_7_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_7_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_7_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_7_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_7_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_7_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_7_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_7_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_7_ARID : IN STD_LOGIC;
    twiddle_rsc_0_7_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_7_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_7_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_7_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_7_BID : OUT STD_LOGIC;
    twiddle_rsc_0_7_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_7_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_7_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_7_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_7_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_7_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_7_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_7_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_7_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_7_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_7_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_7_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_7_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_7_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_7_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_7_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_rsc_0_8_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_8_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_8_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_8_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_8_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_8_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_8_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_8_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_8_RID : OUT STD_LOGIC;
    twiddle_rsc_0_8_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_8_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_8_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_8_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_8_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_8_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_8_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_8_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_8_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_8_ARID : IN STD_LOGIC;
    twiddle_rsc_0_8_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_8_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_8_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_8_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_8_BID : OUT STD_LOGIC;
    twiddle_rsc_0_8_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_8_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_8_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_8_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_8_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_8_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_8_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_8_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_8_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_8_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_8_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_8_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_8_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_8_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_8_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_8_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_rsc_0_9_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_9_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_9_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_9_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_9_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_9_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_9_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_9_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_9_RID : OUT STD_LOGIC;
    twiddle_rsc_0_9_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_9_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_9_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_9_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_9_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_9_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_9_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_9_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_9_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_9_ARID : IN STD_LOGIC;
    twiddle_rsc_0_9_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_9_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_9_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_9_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_9_BID : OUT STD_LOGIC;
    twiddle_rsc_0_9_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_9_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_9_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_9_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_9_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_9_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_9_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_9_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_9_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_9_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_9_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_9_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_9_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_9_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_9_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_9_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_rsc_0_10_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_10_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_10_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_10_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_10_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_10_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_10_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_10_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_10_RID : OUT STD_LOGIC;
    twiddle_rsc_0_10_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_10_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_10_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_10_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_10_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_10_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_10_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_10_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_10_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_10_ARID : IN STD_LOGIC;
    twiddle_rsc_0_10_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_10_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_10_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_10_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_10_BID : OUT STD_LOGIC;
    twiddle_rsc_0_10_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_10_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_10_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_10_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_10_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_10_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_10_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_10_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_10_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_10_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_10_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_10_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_10_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_10_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_10_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_10_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_rsc_0_11_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_11_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_11_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_11_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_11_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_11_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_11_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_11_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_11_RID : OUT STD_LOGIC;
    twiddle_rsc_0_11_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_11_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_11_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_11_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_11_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_11_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_11_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_11_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_11_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_11_ARID : IN STD_LOGIC;
    twiddle_rsc_0_11_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_11_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_11_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_11_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_11_BID : OUT STD_LOGIC;
    twiddle_rsc_0_11_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_11_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_11_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_11_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_11_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_11_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_11_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_11_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_11_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_11_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_11_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_11_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_11_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_11_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_11_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_11_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_rsc_0_12_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_12_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_12_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_12_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_12_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_12_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_12_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_12_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_12_RID : OUT STD_LOGIC;
    twiddle_rsc_0_12_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_12_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_12_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_12_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_12_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_12_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_12_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_12_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_12_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_12_ARID : IN STD_LOGIC;
    twiddle_rsc_0_12_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_12_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_12_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_12_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_12_BID : OUT STD_LOGIC;
    twiddle_rsc_0_12_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_12_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_12_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_12_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_12_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_12_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_12_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_12_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_12_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_12_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_12_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_12_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_12_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_12_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_12_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_12_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_rsc_0_13_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_13_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_13_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_13_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_13_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_13_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_13_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_13_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_13_RID : OUT STD_LOGIC;
    twiddle_rsc_0_13_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_13_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_13_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_13_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_13_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_13_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_13_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_13_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_13_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_13_ARID : IN STD_LOGIC;
    twiddle_rsc_0_13_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_13_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_13_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_13_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_13_BID : OUT STD_LOGIC;
    twiddle_rsc_0_13_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_13_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_13_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_13_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_13_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_13_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_13_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_13_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_13_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_13_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_13_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_13_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_13_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_13_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_13_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_13_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_rsc_0_14_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_14_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_14_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_14_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_14_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_14_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_14_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_14_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_14_RID : OUT STD_LOGIC;
    twiddle_rsc_0_14_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_14_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_14_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_14_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_14_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_14_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_14_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_14_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_14_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_14_ARID : IN STD_LOGIC;
    twiddle_rsc_0_14_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_14_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_14_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_14_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_14_BID : OUT STD_LOGIC;
    twiddle_rsc_0_14_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_14_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_14_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_14_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_14_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_14_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_14_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_14_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_14_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_14_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_14_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_14_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_14_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_14_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_14_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_14_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_rsc_0_15_s_tdone : IN STD_LOGIC;
    twiddle_rsc_0_15_tr_write_done : IN STD_LOGIC;
    twiddle_rsc_0_15_RREADY : IN STD_LOGIC;
    twiddle_rsc_0_15_RVALID : OUT STD_LOGIC;
    twiddle_rsc_0_15_RUSER : OUT STD_LOGIC;
    twiddle_rsc_0_15_RLAST : OUT STD_LOGIC;
    twiddle_rsc_0_15_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_15_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_15_RID : OUT STD_LOGIC;
    twiddle_rsc_0_15_ARREADY : OUT STD_LOGIC;
    twiddle_rsc_0_15_ARVALID : IN STD_LOGIC;
    twiddle_rsc_0_15_ARUSER : IN STD_LOGIC;
    twiddle_rsc_0_15_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_15_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_ARLOCK : IN STD_LOGIC;
    twiddle_rsc_0_15_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_15_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_15_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_15_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_15_ARID : IN STD_LOGIC;
    twiddle_rsc_0_15_BREADY : IN STD_LOGIC;
    twiddle_rsc_0_15_BVALID : OUT STD_LOGIC;
    twiddle_rsc_0_15_BUSER : OUT STD_LOGIC;
    twiddle_rsc_0_15_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_15_BID : OUT STD_LOGIC;
    twiddle_rsc_0_15_WREADY : OUT STD_LOGIC;
    twiddle_rsc_0_15_WVALID : IN STD_LOGIC;
    twiddle_rsc_0_15_WUSER : IN STD_LOGIC;
    twiddle_rsc_0_15_WLAST : IN STD_LOGIC;
    twiddle_rsc_0_15_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_rsc_0_15_AWREADY : OUT STD_LOGIC;
    twiddle_rsc_0_15_AWVALID : IN STD_LOGIC;
    twiddle_rsc_0_15_AWUSER : IN STD_LOGIC;
    twiddle_rsc_0_15_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_15_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_rsc_0_15_AWLOCK : IN STD_LOGIC;
    twiddle_rsc_0_15_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_rsc_0_15_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_rsc_0_15_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_rsc_0_15_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_rsc_0_15_AWID : IN STD_LOGIC;
    twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_0_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_0_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_0_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_0_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_0_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_0_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_0_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_0_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_0_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_0_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_0_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_0_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_0_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_0_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_0_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_1_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_1_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_1_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_1_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_1_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_1_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_1_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_1_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_1_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_1_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_1_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_1_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_1_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_1_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_1_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_1_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_1_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_1_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_1_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_1_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_1_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_1_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_1_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_1_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_1_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_1_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_1_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_1_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_1_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_2_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_2_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_2_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_2_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_2_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_2_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_2_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_2_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_2_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_2_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_2_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_2_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_2_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_2_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_2_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_2_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_2_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_2_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_2_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_2_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_2_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_2_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_2_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_2_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_2_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_2_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_2_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_2_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_2_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_3_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_3_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_3_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_3_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_3_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_3_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_3_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_3_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_3_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_3_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_3_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_3_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_3_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_3_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_3_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_3_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_3_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_3_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_3_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_3_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_3_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_3_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_3_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_3_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_3_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_3_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_3_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_3_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_3_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_4_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_4_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_4_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_4_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_4_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_4_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_4_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_4_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_4_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_4_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_4_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_4_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_4_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_4_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_4_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_4_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_4_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_4_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_4_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_4_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_4_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_4_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_4_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_4_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_4_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_4_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_4_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_4_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_4_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_5_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_5_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_5_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_5_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_5_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_5_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_5_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_5_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_5_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_5_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_5_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_5_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_5_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_5_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_5_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_5_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_5_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_5_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_5_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_5_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_5_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_5_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_5_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_5_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_5_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_5_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_5_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_5_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_5_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_6_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_6_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_6_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_6_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_6_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_6_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_6_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_6_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_6_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_6_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_6_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_6_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_6_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_6_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_6_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_6_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_6_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_6_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_6_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_6_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_6_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_6_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_6_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_6_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_6_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_6_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_6_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_6_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_6_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_7_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_7_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_7_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_7_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_7_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_7_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_7_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_7_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_7_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_7_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_7_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_7_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_7_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_7_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_7_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_7_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_7_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_7_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_7_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_7_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_7_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_7_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_7_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_7_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_7_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_7_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_7_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_7_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_7_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_8_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_8_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_8_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_8_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_8_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_8_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_8_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_8_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_8_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_8_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_8_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_8_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_8_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_8_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_8_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_8_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_8_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_8_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_8_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_8_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_8_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_8_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_8_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_8_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_8_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_8_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_8_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_8_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_8_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_8_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_8_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_9_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_9_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_9_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_9_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_9_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_9_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_9_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_9_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_9_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_9_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_9_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_9_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_9_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_9_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_9_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_9_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_9_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_9_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_9_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_9_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_9_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_9_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_9_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_9_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_9_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_9_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_9_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_9_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_9_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_9_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_9_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_10_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_10_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_10_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_10_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_10_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_10_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_10_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_10_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_10_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_10_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_10_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_10_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_10_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_10_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_10_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_10_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_10_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_10_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_10_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_10_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_10_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_10_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_10_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_10_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_10_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_10_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_10_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_10_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_10_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_10_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_10_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_11_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_11_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_11_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_11_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_11_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_11_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_11_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_11_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_11_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_11_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_11_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_11_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_11_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_11_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_11_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_11_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_11_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_11_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_11_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_11_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_11_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_11_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_11_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_11_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_11_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_11_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_11_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_11_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_11_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_11_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_11_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_12_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_12_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_12_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_12_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_12_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_12_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_12_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_12_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_12_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_12_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_12_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_12_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_12_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_12_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_12_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_12_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_12_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_12_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_12_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_12_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_12_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_12_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_12_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_12_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_12_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_12_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_12_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_12_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_12_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_12_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_12_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_13_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_13_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_13_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_13_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_13_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_13_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_13_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_13_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_13_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_13_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_13_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_13_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_13_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_13_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_13_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_13_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_13_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_13_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_13_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_13_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_13_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_13_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_13_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_13_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_13_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_13_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_13_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_13_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_13_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_13_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_13_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_14_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_14_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_14_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_14_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_14_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_14_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_14_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_14_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_14_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_14_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_14_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_14_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_14_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_14_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_14_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_14_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_14_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_14_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_14_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_14_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_14_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_14_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_14_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_14_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_14_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_14_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_14_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_14_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_14_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_14_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_14_lz : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_s_tdone : IN STD_LOGIC;
    twiddle_h_rsc_0_15_tr_write_done : IN STD_LOGIC;
    twiddle_h_rsc_0_15_RREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_15_RVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_RUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_RLAST : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_15_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_15_RID : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_ARREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_ARVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_15_ARUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_15_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_15_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_ARLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_15_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_15_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_15_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_15_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_15_ARID : IN STD_LOGIC;
    twiddle_h_rsc_0_15_BREADY : IN STD_LOGIC;
    twiddle_h_rsc_0_15_BVALID : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_BUSER : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_15_BID : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_WREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_WVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_15_WUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_15_WLAST : IN STD_LOGIC;
    twiddle_h_rsc_0_15_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
    twiddle_h_rsc_0_15_AWREADY : OUT STD_LOGIC;
    twiddle_h_rsc_0_15_AWVALID : IN STD_LOGIC;
    twiddle_h_rsc_0_15_AWUSER : IN STD_LOGIC;
    twiddle_h_rsc_0_15_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_15_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
    twiddle_h_rsc_0_15_AWLOCK : IN STD_LOGIC;
    twiddle_h_rsc_0_15_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
    twiddle_h_rsc_0_15_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    twiddle_h_rsc_0_15_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
    twiddle_h_rsc_0_15_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    twiddle_h_rsc_0_15_AWID : IN STD_LOGIC;
    twiddle_h_rsc_triosy_0_15_lz : OUT STD_LOGIC
  );
END peaseNTT;

ARCHITECTURE v29 OF peaseNTT IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';
  CONSTANT GND : STD_LOGIC := '0';

  -- Interconnect Declarations
  SIGNAL yt_rsc_0_0_i_clken_d : STD_LOGIC;
  SIGNAL yt_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_clken_d : STD_LOGIC;
  SIGNAL yt_rsc_0_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_clken_d : STD_LOGIC;
  SIGNAL yt_rsc_1_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_clken_d : STD_LOGIC;
  SIGNAL yt_rsc_1_16_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_0_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL xt_rsc_1_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : STD_LOGIC;
  SIGNAL yt_rsc_0_0_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_0_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_1_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_1_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_1_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_2_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_2_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_2_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_3_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_3_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_3_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_4_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_4_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_4_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_5_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_5_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_5_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_6_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_6_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_6_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_7_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_7_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_7_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_8_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_8_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_8_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_9_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_9_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_9_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_10_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_10_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_10_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_11_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_11_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_11_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_12_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_12_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_12_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_13_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_13_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_13_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_14_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_14_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_14_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_15_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_15_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_15_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_16_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_16_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_16_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_17_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_17_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_17_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_18_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_18_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_18_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_19_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_19_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_19_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_20_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_20_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_20_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_21_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_21_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_21_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_22_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_22_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_22_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_23_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_23_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_23_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_24_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_24_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_24_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_25_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_25_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_25_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_26_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_26_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_26_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_27_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_27_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_27_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_28_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_28_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_28_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_29_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_29_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_29_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_30_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_30_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_30_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_clken : STD_LOGIC;
  SIGNAL yt_rsc_0_31_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_wea : STD_LOGIC;
  SIGNAL yt_rsc_0_31_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_31_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_0_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_0_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_0_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_1_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_1_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_1_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_2_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_2_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_2_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_3_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_3_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_3_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_4_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_4_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_4_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_5_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_5_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_5_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_6_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_6_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_6_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_7_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_7_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_7_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_8_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_8_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_8_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_9_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_9_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_9_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_10_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_10_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_10_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_11_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_11_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_11_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_12_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_12_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_12_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_13_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_13_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_13_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_14_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_14_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_14_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_15_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_15_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_15_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_16_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_16_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_16_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_17_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_17_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_17_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_18_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_18_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_18_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_19_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_19_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_19_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_20_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_20_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_20_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_21_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_21_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_21_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_22_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_22_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_22_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_23_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_23_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_23_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_24_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_24_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_24_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_25_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_25_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_25_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_26_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_26_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_26_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_27_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_27_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_27_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_28_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_28_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_28_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_29_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_29_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_29_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_30_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_30_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_30_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_clken : STD_LOGIC;
  SIGNAL yt_rsc_1_31_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_wea : STD_LOGIC;
  SIGNAL yt_rsc_1_31_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_31_unc_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_wea_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_0_1_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_wea_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_1_0_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_wea_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff : STD_LOGIC;
  SIGNAL yt_rsc_1_16_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_0_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_1_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_2_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_3_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_4_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_5_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_6_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_7_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_8_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_9_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_10_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_11_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_12_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_13_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_14_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_15_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_16_i_adra_d_iff : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_17_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_18_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_19_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_20_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_21_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_22_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_23_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_24_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_25_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_26_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_27_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_28_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_29_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_30_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_0_31_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_0_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_0_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_1_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_1_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_2_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_2_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_3_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_3_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_4_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_4_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_5_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_5_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_6_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_6_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_7_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_7_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_8_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_8_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_9_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_9_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_10_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_10_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_11_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_11_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_12_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_12_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_13_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_13_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_14_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_14_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_15_i_da_d_iff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_15_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_16_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_17_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_18_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_19_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_20_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_21_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_22_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_23_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_24_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_25_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_26_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_27_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_28_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_29_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_30_i_wea_d_iff : STD_LOGIC;
  SIGNAL xt_rsc_1_31_i_wea_d_iff : STD_LOGIC;

  SIGNAL yt_rsc_0_0_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_0_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_1_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_1_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_1_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_2_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_2_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_2_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_3_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_3_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_3_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_4_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_4_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_4_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_5_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_5_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_5_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_6_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_6_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_6_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_7_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_7_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_7_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_8_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_8_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_8_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_9_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_9_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_9_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_10_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_10_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_10_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_11_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_11_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_11_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_12_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_12_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_12_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_13_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_13_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_13_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_14_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_14_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_14_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_15_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_15_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_15_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_16_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_16_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_16_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_17_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_17_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_17_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_18_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_18_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_18_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_19_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_19_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_19_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_20_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_20_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_20_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_21_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_21_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_21_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_22_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_22_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_22_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_23_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_23_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_23_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_24_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_24_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_24_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_25_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_25_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_25_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_26_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_26_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_26_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_27_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_27_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_27_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_28_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_28_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_28_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_29_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_29_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_29_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_30_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_30_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_30_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_0_31_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_31_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_31_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_0_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_0_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_0_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_1_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_1_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_1_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_2_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_2_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_2_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_3_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_3_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_3_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_4_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_4_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_4_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_5_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_5_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_5_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_6_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_6_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_6_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_7_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_7_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_7_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_8_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_8_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_8_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_9_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_9_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_9_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_10_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_10_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_10_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_11_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_11_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_11_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_12_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_12_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_12_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_13_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_13_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_13_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_14_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_14_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_14_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_15_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_15_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_15_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_16_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_16_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_16_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_17_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_17_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_17_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_18_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_18_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_18_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_19_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_19_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_19_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_20_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_20_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_20_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_21_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_21_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_21_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_22_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_22_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_22_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_23_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_23_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_23_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_24_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_24_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_24_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_25_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_25_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_25_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_26_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_26_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_26_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_27_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_27_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_27_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_28_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_28_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_28_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_29_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_29_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_29_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_30_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_30_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_30_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  SIGNAL yt_rsc_1_31_comp_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_31_comp_adrb : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_31_comp_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_comp_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_comp_qb : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_7_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_8_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_1_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_9_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_2_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_10_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_3_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_11_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_4_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_12_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_5_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_13_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_6_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_14_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_7_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_15_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_8_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_16_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_9_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_17_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_10_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_18_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_11_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_19_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_12_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_20_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_13_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_21_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_14_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_22_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_15_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_23_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_16_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_16_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_24_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_17_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_17_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_25_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_18_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_18_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_26_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_19_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_19_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_27_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_20_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_20_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_28_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_21_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_21_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_29_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_22_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_22_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_30_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_23_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_23_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_31_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_24_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_24_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_32_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_25_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_25_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_33_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_26_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_26_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_34_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_27_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_27_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_35_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_28_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_28_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_36_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_29_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_29_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_37_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_30_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_30_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_38_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_0_31_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_0_31_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_39_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_0_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_40_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_1_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_41_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_2_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_42_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_3_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_43_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_4_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_44_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_5_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_45_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_6_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_46_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_7_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_47_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_8_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_48_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_9_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_49_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_10_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_50_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_11_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_51_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_12_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_52_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_13_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_53_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_14_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_54_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_15_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_55_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_16_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_16_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_56_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_17_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_17_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_57_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_18_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_18_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_58_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_19_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_19_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_59_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_20_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_20_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_60_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_21_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_21_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_61_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_22_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_22_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_62_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_23_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_23_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_63_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_24_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_24_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_64_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_25_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_25_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_65_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_26_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_26_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_66_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_27_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_27_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_67_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_28_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_28_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_68_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_29_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_29_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_69_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_30_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_30_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_70_4_32_16_16_32_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL yt_rsc_1_31_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_da_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL yt_rsc_1_31_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_71_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_0_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_72_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_1_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_73_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_2_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_74_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_3_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_75_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_4_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_76_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_5_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_77_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_6_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_78_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_7_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_79_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_8_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_80_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_9_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_81_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_10_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_82_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_11_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_83_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_12_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_84_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_13_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_85_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_14_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_86_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_15_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_87_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_16_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_16_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_88_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_17_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_17_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_89_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_18_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_18_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_90_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_19_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_19_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_91_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_20_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_20_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_92_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_21_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_21_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_93_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_22_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_22_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_94_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_23_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_23_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_95_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_24_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_24_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_96_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_25_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_25_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_97_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_26_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_26_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_98_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_27_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_27_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_99_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_28_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_28_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_100_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_29_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_29_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_101_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_30_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_30_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_102_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_0_31_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_0_31_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_103_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_0_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_0_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_0_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_0_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_0_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_104_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_1_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_1_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_1_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_1_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_1_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_105_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_2_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_2_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_2_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_2_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_2_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_106_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_3_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_3_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_3_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_3_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_3_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_107_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_4_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_4_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_4_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_4_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_4_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_108_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_5_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_5_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_5_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_5_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_5_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_109_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_6_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_6_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_6_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_6_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_6_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_110_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_7_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_7_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_7_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_7_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_7_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_111_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_8_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_8_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_8_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_8_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_8_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_8_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_112_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_9_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_9_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_9_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_9_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_9_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_9_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_113_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_10_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_10_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_10_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_10_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_10_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_10_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_114_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_11_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_11_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_11_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_11_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_11_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_11_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_115_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_12_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_12_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_12_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_12_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_12_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_12_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_116_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_13_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_13_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_13_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_13_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_13_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_13_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_117_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_14_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_14_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_14_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_14_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_14_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_14_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_118_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_15_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_15_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_15_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_15_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_15_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_15_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_119_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_16_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_16_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_16_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_16_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_16_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_16_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_120_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_17_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_17_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_17_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_17_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_17_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_17_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_121_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_18_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_18_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_18_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_18_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_18_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_18_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_122_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_19_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_19_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_19_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_19_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_19_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_19_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_123_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_20_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_20_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_20_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_20_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_20_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_20_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_124_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_21_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_21_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_21_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_21_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_21_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_21_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_125_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_22_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_22_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_22_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_22_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_22_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_22_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_126_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_23_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_23_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_23_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_23_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_23_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_23_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_127_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_24_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_24_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_24_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_24_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_24_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_24_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_128_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_25_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_25_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_25_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_25_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_25_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_25_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_129_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_26_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_26_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_26_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_26_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_26_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_26_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_130_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_27_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_27_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_27_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_27_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_27_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_27_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_131_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_28_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_28_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_28_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_28_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_28_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_28_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_132_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_29_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_29_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_29_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_29_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_29_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_29_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_133_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_30_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_30_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_30_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_30_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_30_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_30_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_134_4_32_16_16_32_1_gen
    PORT(
      qa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea : OUT STD_LOGIC;
      da : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      adra : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      adra_d : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      da_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      qa_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      wea_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_RMASK_B_d : IN STD_LOGIC;
      rwA_rw_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL xt_rsc_1_31_i_qa : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_31_i_da : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_31_i_adra : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_31_i_adra_d : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL xt_rsc_1_31_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL xt_rsc_1_31_i_qa_d_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);

  COMPONENT peaseNTT_core
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      xt_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_16_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_17_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_18_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_19_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_20_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_21_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_22_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_23_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_24_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_25_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_26_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_27_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_28_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_29_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_30_lz : OUT STD_LOGIC;
      xt_rsc_triosy_0_31_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_0_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_1_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_2_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_3_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_4_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_5_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_6_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_7_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_8_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_9_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_10_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_11_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_12_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_13_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_14_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_15_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_16_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_17_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_18_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_19_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_20_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_21_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_22_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_23_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_24_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_25_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_26_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_27_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_28_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_29_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_30_lz : OUT STD_LOGIC;
      xt_rsc_triosy_1_31_lz : OUT STD_LOGIC;
      p_rsc_dat : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      p_rsc_triosy_lz : OUT STD_LOGIC;
      r_rsc_triosy_lz : OUT STD_LOGIC;
      twiddle_rsc_0_0_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_0_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_0_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_0_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_0_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_0_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_0_RID : OUT STD_LOGIC;
      twiddle_rsc_0_0_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_0_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_0_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_0_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_0_ARID : IN STD_LOGIC;
      twiddle_rsc_0_0_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_0_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_0_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_0_BID : OUT STD_LOGIC;
      twiddle_rsc_0_0_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_0_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_0_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_0_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_0_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_0_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_0_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_0_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_0_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      twiddle_rsc_0_1_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_1_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_1_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_1_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_1_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_1_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_1_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_1_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_1_RID : OUT STD_LOGIC;
      twiddle_rsc_0_1_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_1_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_1_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_1_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_1_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_1_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_1_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_1_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_1_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_1_ARID : IN STD_LOGIC;
      twiddle_rsc_0_1_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_1_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_1_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_1_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_1_BID : OUT STD_LOGIC;
      twiddle_rsc_0_1_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_1_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_1_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_1_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_1_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_1_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_1_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_1_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_1_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_1_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_1_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_1_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_1_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_1_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_1_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_1_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      twiddle_rsc_0_2_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_2_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_2_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_2_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_2_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_2_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_2_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_2_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_2_RID : OUT STD_LOGIC;
      twiddle_rsc_0_2_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_2_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_2_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_2_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_2_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_2_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_2_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_2_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_2_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_2_ARID : IN STD_LOGIC;
      twiddle_rsc_0_2_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_2_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_2_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_2_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_2_BID : OUT STD_LOGIC;
      twiddle_rsc_0_2_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_2_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_2_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_2_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_2_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_2_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_2_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_2_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_2_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_2_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_2_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_2_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_2_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_2_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_2_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_2_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      twiddle_rsc_0_3_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_3_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_3_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_3_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_3_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_3_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_3_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_3_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_3_RID : OUT STD_LOGIC;
      twiddle_rsc_0_3_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_3_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_3_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_3_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_3_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_3_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_3_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_3_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_3_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_3_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_3_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_3_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_3_ARID : IN STD_LOGIC;
      twiddle_rsc_0_3_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_3_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_3_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_3_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_3_BID : OUT STD_LOGIC;
      twiddle_rsc_0_3_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_3_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_3_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_3_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_3_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_3_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_3_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_3_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_3_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_3_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_3_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_3_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_3_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_3_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_3_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_3_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_3_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_3_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_3_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      twiddle_rsc_0_4_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_4_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_4_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_4_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_4_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_4_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_4_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_4_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_4_RID : OUT STD_LOGIC;
      twiddle_rsc_0_4_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_4_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_4_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_4_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_4_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_4_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_4_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_4_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_4_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_4_ARID : IN STD_LOGIC;
      twiddle_rsc_0_4_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_4_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_4_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_4_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_4_BID : OUT STD_LOGIC;
      twiddle_rsc_0_4_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_4_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_4_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_4_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_4_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_4_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_4_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_4_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_4_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_4_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_4_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_4_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_4_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_4_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_4_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_4_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      twiddle_rsc_0_5_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_5_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_5_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_5_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_5_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_5_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_5_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_5_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_5_RID : OUT STD_LOGIC;
      twiddle_rsc_0_5_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_5_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_5_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_5_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_5_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_5_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_5_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_5_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_5_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_5_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_5_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_5_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_5_ARID : IN STD_LOGIC;
      twiddle_rsc_0_5_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_5_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_5_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_5_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_5_BID : OUT STD_LOGIC;
      twiddle_rsc_0_5_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_5_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_5_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_5_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_5_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_5_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_5_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_5_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_5_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_5_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_5_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_5_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_5_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_5_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_5_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_5_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_5_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_5_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_5_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      twiddle_rsc_0_6_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_6_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_6_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_6_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_6_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_6_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_6_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_6_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_6_RID : OUT STD_LOGIC;
      twiddle_rsc_0_6_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_6_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_6_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_6_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_6_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_6_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_6_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_6_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_6_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_6_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_6_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_6_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_6_ARID : IN STD_LOGIC;
      twiddle_rsc_0_6_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_6_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_6_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_6_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_6_BID : OUT STD_LOGIC;
      twiddle_rsc_0_6_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_6_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_6_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_6_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_6_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_6_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_6_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_6_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_6_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_6_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_6_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_6_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_6_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_6_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_6_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_6_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_6_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_6_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_6_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      twiddle_rsc_0_7_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_7_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_7_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_7_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_7_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_7_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_7_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_7_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_7_RID : OUT STD_LOGIC;
      twiddle_rsc_0_7_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_7_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_7_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_7_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_7_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_7_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_7_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_7_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_7_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_7_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_7_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_7_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_7_ARID : IN STD_LOGIC;
      twiddle_rsc_0_7_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_7_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_7_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_7_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_7_BID : OUT STD_LOGIC;
      twiddle_rsc_0_7_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_7_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_7_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_7_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_7_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_7_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_7_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_7_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_7_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_7_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_7_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_7_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_7_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_7_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_7_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_7_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_7_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_7_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_7_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      twiddle_rsc_0_8_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_8_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_8_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_8_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_8_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_8_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_8_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_8_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_8_RID : OUT STD_LOGIC;
      twiddle_rsc_0_8_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_8_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_8_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_8_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_8_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_8_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_8_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_8_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_8_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_8_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_8_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_8_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_8_ARID : IN STD_LOGIC;
      twiddle_rsc_0_8_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_8_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_8_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_8_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_8_BID : OUT STD_LOGIC;
      twiddle_rsc_0_8_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_8_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_8_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_8_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_8_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_8_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_8_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_8_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_8_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_8_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_8_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_8_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_8_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_8_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_8_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_8_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_8_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_8_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_8_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      twiddle_rsc_0_9_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_9_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_9_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_9_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_9_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_9_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_9_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_9_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_9_RID : OUT STD_LOGIC;
      twiddle_rsc_0_9_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_9_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_9_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_9_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_9_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_9_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_9_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_9_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_9_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_9_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_9_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_9_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_9_ARID : IN STD_LOGIC;
      twiddle_rsc_0_9_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_9_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_9_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_9_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_9_BID : OUT STD_LOGIC;
      twiddle_rsc_0_9_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_9_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_9_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_9_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_9_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_9_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_9_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_9_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_9_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_9_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_9_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_9_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_9_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_9_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_9_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_9_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_9_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_9_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_9_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      twiddle_rsc_0_10_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_10_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_10_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_10_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_10_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_10_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_10_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_10_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_10_RID : OUT STD_LOGIC;
      twiddle_rsc_0_10_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_10_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_10_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_10_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_10_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_10_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_10_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_10_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_10_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_10_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_10_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_10_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_10_ARID : IN STD_LOGIC;
      twiddle_rsc_0_10_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_10_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_10_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_10_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_10_BID : OUT STD_LOGIC;
      twiddle_rsc_0_10_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_10_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_10_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_10_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_10_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_10_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_10_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_10_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_10_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_10_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_10_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_10_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_10_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_10_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_10_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_10_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_10_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_10_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_10_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      twiddle_rsc_0_11_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_11_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_11_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_11_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_11_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_11_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_11_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_11_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_11_RID : OUT STD_LOGIC;
      twiddle_rsc_0_11_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_11_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_11_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_11_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_11_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_11_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_11_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_11_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_11_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_11_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_11_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_11_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_11_ARID : IN STD_LOGIC;
      twiddle_rsc_0_11_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_11_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_11_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_11_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_11_BID : OUT STD_LOGIC;
      twiddle_rsc_0_11_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_11_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_11_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_11_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_11_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_11_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_11_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_11_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_11_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_11_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_11_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_11_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_11_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_11_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_11_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_11_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_11_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_11_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_11_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      twiddle_rsc_0_12_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_12_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_12_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_12_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_12_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_12_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_12_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_12_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_12_RID : OUT STD_LOGIC;
      twiddle_rsc_0_12_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_12_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_12_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_12_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_12_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_12_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_12_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_12_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_12_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_12_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_12_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_12_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_12_ARID : IN STD_LOGIC;
      twiddle_rsc_0_12_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_12_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_12_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_12_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_12_BID : OUT STD_LOGIC;
      twiddle_rsc_0_12_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_12_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_12_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_12_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_12_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_12_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_12_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_12_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_12_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_12_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_12_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_12_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_12_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_12_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_12_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_12_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_12_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_12_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_12_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      twiddle_rsc_0_13_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_13_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_13_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_13_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_13_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_13_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_13_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_13_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_13_RID : OUT STD_LOGIC;
      twiddle_rsc_0_13_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_13_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_13_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_13_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_13_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_13_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_13_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_13_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_13_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_13_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_13_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_13_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_13_ARID : IN STD_LOGIC;
      twiddle_rsc_0_13_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_13_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_13_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_13_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_13_BID : OUT STD_LOGIC;
      twiddle_rsc_0_13_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_13_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_13_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_13_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_13_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_13_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_13_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_13_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_13_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_13_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_13_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_13_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_13_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_13_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_13_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_13_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_13_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_13_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_13_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      twiddle_rsc_0_14_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_14_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_14_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_14_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_14_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_14_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_14_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_14_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_14_RID : OUT STD_LOGIC;
      twiddle_rsc_0_14_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_14_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_14_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_14_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_14_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_14_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_14_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_14_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_14_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_14_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_14_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_14_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_14_ARID : IN STD_LOGIC;
      twiddle_rsc_0_14_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_14_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_14_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_14_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_14_BID : OUT STD_LOGIC;
      twiddle_rsc_0_14_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_14_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_14_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_14_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_14_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_14_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_14_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_14_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_14_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_14_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_14_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_14_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_14_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_14_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_14_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_14_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_14_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_14_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_14_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      twiddle_rsc_0_15_s_tdone : IN STD_LOGIC;
      twiddle_rsc_0_15_tr_write_done : IN STD_LOGIC;
      twiddle_rsc_0_15_RREADY : IN STD_LOGIC;
      twiddle_rsc_0_15_RVALID : OUT STD_LOGIC;
      twiddle_rsc_0_15_RUSER : OUT STD_LOGIC;
      twiddle_rsc_0_15_RLAST : OUT STD_LOGIC;
      twiddle_rsc_0_15_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_15_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_15_RID : OUT STD_LOGIC;
      twiddle_rsc_0_15_ARREADY : OUT STD_LOGIC;
      twiddle_rsc_0_15_ARVALID : IN STD_LOGIC;
      twiddle_rsc_0_15_ARUSER : IN STD_LOGIC;
      twiddle_rsc_0_15_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_15_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_15_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_15_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_15_ARLOCK : IN STD_LOGIC;
      twiddle_rsc_0_15_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_15_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_15_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_15_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_15_ARID : IN STD_LOGIC;
      twiddle_rsc_0_15_BREADY : IN STD_LOGIC;
      twiddle_rsc_0_15_BVALID : OUT STD_LOGIC;
      twiddle_rsc_0_15_BUSER : OUT STD_LOGIC;
      twiddle_rsc_0_15_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_15_BID : OUT STD_LOGIC;
      twiddle_rsc_0_15_WREADY : OUT STD_LOGIC;
      twiddle_rsc_0_15_WVALID : IN STD_LOGIC;
      twiddle_rsc_0_15_WUSER : IN STD_LOGIC;
      twiddle_rsc_0_15_WLAST : IN STD_LOGIC;
      twiddle_rsc_0_15_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_15_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_rsc_0_15_AWREADY : OUT STD_LOGIC;
      twiddle_rsc_0_15_AWVALID : IN STD_LOGIC;
      twiddle_rsc_0_15_AWUSER : IN STD_LOGIC;
      twiddle_rsc_0_15_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_15_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_15_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_15_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_rsc_0_15_AWLOCK : IN STD_LOGIC;
      twiddle_rsc_0_15_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_rsc_0_15_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_rsc_0_15_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_rsc_0_15_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_rsc_0_15_AWID : IN STD_LOGIC;
      twiddle_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_0_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_0_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_0_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_0_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_0_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_0_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_0_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_0_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_0_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_0_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_0_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_0_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_0_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_0_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_0_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_0_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_0_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_0_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_0_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_0_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_0_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_0_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_0_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_0_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_0_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_0_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_0_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_0_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_0_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_0_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_0_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_0_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_0_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_0_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_0_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_0_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_0_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_1_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_1_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_1_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_1_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_1_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_1_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_1_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_1_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_1_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_1_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_1_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_1_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_1_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_1_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_1_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_1_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_1_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_1_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_1_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_1_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_1_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_1_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_1_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_1_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_1_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_1_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_1_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_1_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_1_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_1_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_1_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_1_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_1_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_1_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_1_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_1_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_1_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_2_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_2_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_2_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_2_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_2_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_2_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_2_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_2_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_2_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_2_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_2_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_2_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_2_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_2_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_2_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_2_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_2_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_2_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_2_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_2_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_2_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_2_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_2_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_2_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_2_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_2_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_2_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_2_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_2_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_2_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_2_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_2_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_2_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_2_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_2_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_2_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_2_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_3_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_3_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_3_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_3_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_3_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_3_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_3_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_3_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_3_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_3_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_3_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_3_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_3_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_3_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_3_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_3_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_3_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_3_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_3_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_3_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_3_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_3_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_3_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_3_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_3_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_3_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_3_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_3_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_3_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_3_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_3_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_3_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_3_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_3_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_3_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_3_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_3_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_4_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_4_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_4_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_4_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_4_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_4_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_4_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_4_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_4_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_4_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_4_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_4_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_4_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_4_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_4_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_4_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_4_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_4_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_4_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_4_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_4_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_4_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_4_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_4_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_4_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_4_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_4_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_4_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_4_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_4_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_4_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_4_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_4_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_4_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_4_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_4_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_4_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_5_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_5_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_5_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_5_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_5_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_5_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_5_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_5_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_5_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_5_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_5_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_5_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_5_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_5_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_5_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_5_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_5_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_5_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_5_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_5_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_5_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_5_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_5_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_5_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_5_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_5_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_5_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_5_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_5_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_5_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_5_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_5_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_5_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_5_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_5_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_5_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_5_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_6_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_6_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_6_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_6_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_6_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_6_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_6_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_6_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_6_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_6_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_6_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_6_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_6_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_6_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_6_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_6_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_6_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_6_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_6_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_6_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_6_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_6_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_6_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_6_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_6_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_6_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_6_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_6_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_6_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_6_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_6_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_6_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_6_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_6_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_6_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_6_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_6_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_7_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_7_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_7_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_7_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_7_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_7_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_7_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_7_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_7_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_7_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_7_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_7_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_7_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_7_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_7_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_7_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_7_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_7_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_7_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_7_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_7_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_7_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_7_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_7_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_7_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_7_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_7_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_7_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_7_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_7_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_7_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_7_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_7_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_7_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_7_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_7_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_7_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_8_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_8_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_8_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_8_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_8_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_8_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_8_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_8_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_8_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_8_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_8_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_8_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_8_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_8_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_8_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_8_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_8_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_8_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_8_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_8_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_8_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_8_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_8_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_8_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_8_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_8_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_8_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_8_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_8_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_8_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_8_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_8_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_8_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_8_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_8_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_8_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_8_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_9_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_9_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_9_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_9_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_9_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_9_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_9_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_9_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_9_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_9_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_9_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_9_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_9_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_9_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_9_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_9_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_9_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_9_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_9_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_9_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_9_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_9_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_9_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_9_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_9_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_9_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_9_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_9_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_9_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_9_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_9_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_9_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_9_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_9_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_9_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_9_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_9_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_10_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_10_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_10_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_10_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_10_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_10_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_10_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_10_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_10_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_10_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_10_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_10_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_10_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_10_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_10_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_10_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_10_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_10_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_10_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_10_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_10_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_10_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_10_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_10_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_10_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_10_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_10_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_10_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_10_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_10_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_10_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_10_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_10_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_10_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_10_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_10_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_10_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_11_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_11_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_11_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_11_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_11_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_11_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_11_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_11_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_11_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_11_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_11_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_11_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_11_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_11_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_11_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_11_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_11_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_11_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_11_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_11_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_11_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_11_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_11_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_11_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_11_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_11_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_11_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_11_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_11_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_11_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_11_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_11_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_11_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_11_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_11_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_11_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_11_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_12_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_12_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_12_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_12_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_12_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_12_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_12_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_12_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_12_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_12_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_12_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_12_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_12_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_12_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_12_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_12_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_12_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_12_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_12_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_12_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_12_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_12_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_12_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_12_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_12_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_12_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_12_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_12_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_12_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_12_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_12_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_12_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_12_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_12_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_12_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_12_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_12_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_13_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_13_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_13_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_13_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_13_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_13_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_13_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_13_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_13_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_13_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_13_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_13_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_13_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_13_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_13_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_13_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_13_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_13_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_13_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_13_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_13_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_13_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_13_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_13_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_13_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_13_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_13_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_13_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_13_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_13_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_13_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_13_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_13_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_13_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_13_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_13_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_13_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_14_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_14_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_14_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_14_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_14_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_14_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_14_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_14_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_14_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_14_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_14_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_14_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_14_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_14_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_14_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_14_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_14_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_14_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_14_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_14_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_14_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_14_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_14_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_14_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_14_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_14_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_14_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_14_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_14_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_14_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_14_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_14_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_14_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_14_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_14_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_14_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_14_lz : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_s_tdone : IN STD_LOGIC;
      twiddle_h_rsc_0_15_tr_write_done : IN STD_LOGIC;
      twiddle_h_rsc_0_15_RREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_15_RVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_RUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_RLAST : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_RRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_15_RDATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_15_RID : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_ARREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_ARVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_15_ARUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_15_ARREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_15_ARQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_15_ARPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_15_ARCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_15_ARLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_15_ARBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_15_ARSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_15_ARLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_15_ARADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_15_ARID : IN STD_LOGIC;
      twiddle_h_rsc_0_15_BREADY : IN STD_LOGIC;
      twiddle_h_rsc_0_15_BVALID : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_BUSER : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_BRESP : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_15_BID : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_WREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_WVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_15_WUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_15_WLAST : IN STD_LOGIC;
      twiddle_h_rsc_0_15_WSTRB : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_15_WDATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      twiddle_h_rsc_0_15_AWREADY : OUT STD_LOGIC;
      twiddle_h_rsc_0_15_AWVALID : IN STD_LOGIC;
      twiddle_h_rsc_0_15_AWUSER : IN STD_LOGIC;
      twiddle_h_rsc_0_15_AWREGION : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_15_AWQOS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_15_AWPROT : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_15_AWCACHE : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
      twiddle_h_rsc_0_15_AWLOCK : IN STD_LOGIC;
      twiddle_h_rsc_0_15_AWBURST : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
      twiddle_h_rsc_0_15_AWSIZE : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      twiddle_h_rsc_0_15_AWLEN : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
      twiddle_h_rsc_0_15_AWADDR : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      twiddle_h_rsc_0_15_AWID : IN STD_LOGIC;
      twiddle_h_rsc_triosy_0_15_lz : OUT STD_LOGIC;
      yt_rsc_0_0_i_clken_d : OUT STD_LOGIC;
      yt_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_16_i_clken_d : OUT STD_LOGIC;
      yt_rsc_0_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_0_i_clken_d : OUT STD_LOGIC;
      yt_rsc_1_0_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_1_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_2_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_3_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_4_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_5_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_6_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_7_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_8_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_9_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_10_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_11_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_12_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_13_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_14_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_15_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_16_i_clken_d : OUT STD_LOGIC;
      yt_rsc_1_16_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_17_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_18_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_19_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_20_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_21_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_22_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_23_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_24_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_25_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_26_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_27_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_28_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_29_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_30_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_31_i_da_d : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_1_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_0_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_0_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_1_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_2_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_3_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_4_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_5_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_6_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_7_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_8_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_9_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_10_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_11_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_12_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_13_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_14_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_15_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_16_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_17_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_18_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_19_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_20_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_21_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_22_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_23_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_24_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_25_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_26_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_27_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_28_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_29_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_30_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      xt_rsc_1_31_i_qa_d : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d : OUT STD_LOGIC;
      yt_rsc_0_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
      yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      yt_rsc_0_1_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_2_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_3_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_4_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_5_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_6_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_7_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_8_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_9_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_10_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_11_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_12_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_13_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_14_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_15_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      yt_rsc_0_16_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_0_16_i_wea_d_pff : OUT STD_LOGIC;
      yt_rsc_1_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_1_0_i_wea_d_pff : OUT STD_LOGIC;
      yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff : OUT STD_LOGIC;
      yt_rsc_1_16_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      yt_rsc_1_16_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_0_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_0_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_1_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_1_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_2_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_2_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_3_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_3_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_4_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_4_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_5_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_5_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_6_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_6_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_7_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_7_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_8_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_8_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_9_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_9_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_10_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_10_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_11_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_11_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_12_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_12_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_13_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_13_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_14_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_14_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_15_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_0_15_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_16_i_adra_d_pff : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
      xt_rsc_0_16_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_17_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_18_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_19_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_20_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_21_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_22_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_23_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_24_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_25_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_26_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_27_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_28_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_29_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_30_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_0_31_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_0_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_0_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_1_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_1_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_2_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_2_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_3_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_3_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_4_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_4_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_5_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_5_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_6_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_6_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_7_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_7_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_8_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_8_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_9_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_9_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_10_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_10_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_11_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_11_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_12_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_12_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_13_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_13_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_14_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_14_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_15_i_da_d_pff : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
      xt_rsc_1_15_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_16_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_17_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_18_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_19_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_20_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_21_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_22_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_23_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_24_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_25_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_26_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_27_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_28_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_29_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_30_i_wea_d_pff : OUT STD_LOGIC;
      xt_rsc_1_31_i_wea_d_pff : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL peaseNTT_core_inst_p_rsc_dat : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_1_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_2_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_3_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_4_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_5_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_6_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_7_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_8_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_RDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_WDATA : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_9_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_10_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_11_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_12_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_13_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_14_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_RRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_BRESP : STD_LOGIC_VECTOR (1 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_twiddle_rsc_0_15_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_0_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_1_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_2_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_3_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_4_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_5_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_6_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_7_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_8_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_9_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_10_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_11_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_12_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_13_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_14_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_RRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_RDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_ARREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_ARQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_ARPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_ARCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_ARBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_ARSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_ARLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_ARADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_BRESP : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_WSTRB : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_WDATA : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_AWREGION : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_AWQOS : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_AWPROT : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_AWCACHE : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_AWBURST : STD_LOGIC_VECTOR (1 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_AWSIZE : STD_LOGIC_VECTOR (2 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_AWLEN : STD_LOGIC_VECTOR (7 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_twiddle_h_rsc_0_15_AWADDR : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_0_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_1_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_2_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_3_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_4_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_5_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_6_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_7_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_8_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_9_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_10_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_11_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_12_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_13_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_14_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_15_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_16_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_17_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_18_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_19_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_20_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_21_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_22_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_23_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_24_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_25_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_26_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_27_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_28_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_29_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_30_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_31_i_da_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_0_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_1_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_2_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_3_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_4_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_5_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_6_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_7_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_8_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_9_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_10_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_11_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_12_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_13_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_14_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_15_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_16_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_17_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_18_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_19_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_20_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_21_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_22_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_23_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_24_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_25_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_26_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_27_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_28_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_29_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_30_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_31_i_qa_d : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_0_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_0_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_1_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_2_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_3_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_4_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_5_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_6_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_7_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_8_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_9_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_10_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_11_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_12_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_13_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_14_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_15_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_0_16_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_0_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_yt_rsc_1_16_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_0_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_0_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_1_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_2_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_3_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_4_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_5_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_6_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_7_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_8_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_9_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_10_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_11_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_12_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_13_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_14_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_15_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_0_16_i_adra_d_pff : STD_LOGIC_VECTOR (3 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_0_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_1_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_2_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_3_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_4_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_5_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_6_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_7_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_8_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_9_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO 0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_10_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_11_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_12_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_13_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_14_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);
  SIGNAL peaseNTT_core_inst_xt_rsc_1_15_i_da_d_pff : STD_LOGIC_VECTOR (31 DOWNTO
      0);

BEGIN
  yt_rsc_0_0_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_0_comp_adra,
      adrb => yt_rsc_0_0_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_0_clken,
      da => yt_rsc_0_0_comp_da,
      qa => yt_rsc_0_0_comp_qa,
      qb => yt_rsc_0_0_comp_qb,
      wea => yt_rsc_0_0_wea
    );
  yt_rsc_0_0_comp_adra <= yt_rsc_0_0_adra;
  yt_rsc_0_0_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_0_comp_da <= yt_rsc_0_0_da;
  yt_rsc_0_0_qa <= yt_rsc_0_0_comp_qa;
  yt_rsc_0_0_unc_1 <= yt_rsc_0_0_comp_qb;

  yt_rsc_0_1_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_1_comp_adra,
      adrb => yt_rsc_0_1_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_1_clken,
      da => yt_rsc_0_1_comp_da,
      qa => yt_rsc_0_1_comp_qa,
      qb => yt_rsc_0_1_comp_qb,
      wea => yt_rsc_0_1_wea
    );
  yt_rsc_0_1_comp_adra <= yt_rsc_0_1_adra;
  yt_rsc_0_1_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_1_comp_da <= yt_rsc_0_1_da;
  yt_rsc_0_1_qa <= yt_rsc_0_1_comp_qa;
  yt_rsc_0_1_unc_1 <= yt_rsc_0_1_comp_qb;

  yt_rsc_0_2_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_2_comp_adra,
      adrb => yt_rsc_0_2_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_2_clken,
      da => yt_rsc_0_2_comp_da,
      qa => yt_rsc_0_2_comp_qa,
      qb => yt_rsc_0_2_comp_qb,
      wea => yt_rsc_0_2_wea
    );
  yt_rsc_0_2_comp_adra <= yt_rsc_0_2_adra;
  yt_rsc_0_2_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_2_comp_da <= yt_rsc_0_2_da;
  yt_rsc_0_2_qa <= yt_rsc_0_2_comp_qa;
  yt_rsc_0_2_unc_1 <= yt_rsc_0_2_comp_qb;

  yt_rsc_0_3_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_3_comp_adra,
      adrb => yt_rsc_0_3_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_3_clken,
      da => yt_rsc_0_3_comp_da,
      qa => yt_rsc_0_3_comp_qa,
      qb => yt_rsc_0_3_comp_qb,
      wea => yt_rsc_0_3_wea
    );
  yt_rsc_0_3_comp_adra <= yt_rsc_0_3_adra;
  yt_rsc_0_3_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_3_comp_da <= yt_rsc_0_3_da;
  yt_rsc_0_3_qa <= yt_rsc_0_3_comp_qa;
  yt_rsc_0_3_unc_1 <= yt_rsc_0_3_comp_qb;

  yt_rsc_0_4_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_4_comp_adra,
      adrb => yt_rsc_0_4_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_4_clken,
      da => yt_rsc_0_4_comp_da,
      qa => yt_rsc_0_4_comp_qa,
      qb => yt_rsc_0_4_comp_qb,
      wea => yt_rsc_0_4_wea
    );
  yt_rsc_0_4_comp_adra <= yt_rsc_0_4_adra;
  yt_rsc_0_4_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_4_comp_da <= yt_rsc_0_4_da;
  yt_rsc_0_4_qa <= yt_rsc_0_4_comp_qa;
  yt_rsc_0_4_unc_1 <= yt_rsc_0_4_comp_qb;

  yt_rsc_0_5_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_5_comp_adra,
      adrb => yt_rsc_0_5_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_5_clken,
      da => yt_rsc_0_5_comp_da,
      qa => yt_rsc_0_5_comp_qa,
      qb => yt_rsc_0_5_comp_qb,
      wea => yt_rsc_0_5_wea
    );
  yt_rsc_0_5_comp_adra <= yt_rsc_0_5_adra;
  yt_rsc_0_5_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_5_comp_da <= yt_rsc_0_5_da;
  yt_rsc_0_5_qa <= yt_rsc_0_5_comp_qa;
  yt_rsc_0_5_unc_1 <= yt_rsc_0_5_comp_qb;

  yt_rsc_0_6_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_6_comp_adra,
      adrb => yt_rsc_0_6_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_6_clken,
      da => yt_rsc_0_6_comp_da,
      qa => yt_rsc_0_6_comp_qa,
      qb => yt_rsc_0_6_comp_qb,
      wea => yt_rsc_0_6_wea
    );
  yt_rsc_0_6_comp_adra <= yt_rsc_0_6_adra;
  yt_rsc_0_6_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_6_comp_da <= yt_rsc_0_6_da;
  yt_rsc_0_6_qa <= yt_rsc_0_6_comp_qa;
  yt_rsc_0_6_unc_1 <= yt_rsc_0_6_comp_qb;

  yt_rsc_0_7_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_7_comp_adra,
      adrb => yt_rsc_0_7_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_7_clken,
      da => yt_rsc_0_7_comp_da,
      qa => yt_rsc_0_7_comp_qa,
      qb => yt_rsc_0_7_comp_qb,
      wea => yt_rsc_0_7_wea
    );
  yt_rsc_0_7_comp_adra <= yt_rsc_0_7_adra;
  yt_rsc_0_7_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_7_comp_da <= yt_rsc_0_7_da;
  yt_rsc_0_7_qa <= yt_rsc_0_7_comp_qa;
  yt_rsc_0_7_unc_1 <= yt_rsc_0_7_comp_qb;

  yt_rsc_0_8_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_8_comp_adra,
      adrb => yt_rsc_0_8_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_8_clken,
      da => yt_rsc_0_8_comp_da,
      qa => yt_rsc_0_8_comp_qa,
      qb => yt_rsc_0_8_comp_qb,
      wea => yt_rsc_0_8_wea
    );
  yt_rsc_0_8_comp_adra <= yt_rsc_0_8_adra;
  yt_rsc_0_8_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_8_comp_da <= yt_rsc_0_8_da;
  yt_rsc_0_8_qa <= yt_rsc_0_8_comp_qa;
  yt_rsc_0_8_unc_1 <= yt_rsc_0_8_comp_qb;

  yt_rsc_0_9_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_9_comp_adra,
      adrb => yt_rsc_0_9_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_9_clken,
      da => yt_rsc_0_9_comp_da,
      qa => yt_rsc_0_9_comp_qa,
      qb => yt_rsc_0_9_comp_qb,
      wea => yt_rsc_0_9_wea
    );
  yt_rsc_0_9_comp_adra <= yt_rsc_0_9_adra;
  yt_rsc_0_9_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_9_comp_da <= yt_rsc_0_9_da;
  yt_rsc_0_9_qa <= yt_rsc_0_9_comp_qa;
  yt_rsc_0_9_unc_1 <= yt_rsc_0_9_comp_qb;

  yt_rsc_0_10_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_10_comp_adra,
      adrb => yt_rsc_0_10_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_10_clken,
      da => yt_rsc_0_10_comp_da,
      qa => yt_rsc_0_10_comp_qa,
      qb => yt_rsc_0_10_comp_qb,
      wea => yt_rsc_0_10_wea
    );
  yt_rsc_0_10_comp_adra <= yt_rsc_0_10_adra;
  yt_rsc_0_10_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_10_comp_da <= yt_rsc_0_10_da;
  yt_rsc_0_10_qa <= yt_rsc_0_10_comp_qa;
  yt_rsc_0_10_unc_1 <= yt_rsc_0_10_comp_qb;

  yt_rsc_0_11_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_11_comp_adra,
      adrb => yt_rsc_0_11_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_11_clken,
      da => yt_rsc_0_11_comp_da,
      qa => yt_rsc_0_11_comp_qa,
      qb => yt_rsc_0_11_comp_qb,
      wea => yt_rsc_0_11_wea
    );
  yt_rsc_0_11_comp_adra <= yt_rsc_0_11_adra;
  yt_rsc_0_11_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_11_comp_da <= yt_rsc_0_11_da;
  yt_rsc_0_11_qa <= yt_rsc_0_11_comp_qa;
  yt_rsc_0_11_unc_1 <= yt_rsc_0_11_comp_qb;

  yt_rsc_0_12_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_12_comp_adra,
      adrb => yt_rsc_0_12_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_12_clken,
      da => yt_rsc_0_12_comp_da,
      qa => yt_rsc_0_12_comp_qa,
      qb => yt_rsc_0_12_comp_qb,
      wea => yt_rsc_0_12_wea
    );
  yt_rsc_0_12_comp_adra <= yt_rsc_0_12_adra;
  yt_rsc_0_12_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_12_comp_da <= yt_rsc_0_12_da;
  yt_rsc_0_12_qa <= yt_rsc_0_12_comp_qa;
  yt_rsc_0_12_unc_1 <= yt_rsc_0_12_comp_qb;

  yt_rsc_0_13_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_13_comp_adra,
      adrb => yt_rsc_0_13_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_13_clken,
      da => yt_rsc_0_13_comp_da,
      qa => yt_rsc_0_13_comp_qa,
      qb => yt_rsc_0_13_comp_qb,
      wea => yt_rsc_0_13_wea
    );
  yt_rsc_0_13_comp_adra <= yt_rsc_0_13_adra;
  yt_rsc_0_13_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_13_comp_da <= yt_rsc_0_13_da;
  yt_rsc_0_13_qa <= yt_rsc_0_13_comp_qa;
  yt_rsc_0_13_unc_1 <= yt_rsc_0_13_comp_qb;

  yt_rsc_0_14_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_14_comp_adra,
      adrb => yt_rsc_0_14_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_14_clken,
      da => yt_rsc_0_14_comp_da,
      qa => yt_rsc_0_14_comp_qa,
      qb => yt_rsc_0_14_comp_qb,
      wea => yt_rsc_0_14_wea
    );
  yt_rsc_0_14_comp_adra <= yt_rsc_0_14_adra;
  yt_rsc_0_14_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_14_comp_da <= yt_rsc_0_14_da;
  yt_rsc_0_14_qa <= yt_rsc_0_14_comp_qa;
  yt_rsc_0_14_unc_1 <= yt_rsc_0_14_comp_qb;

  yt_rsc_0_15_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_15_comp_adra,
      adrb => yt_rsc_0_15_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_15_clken,
      da => yt_rsc_0_15_comp_da,
      qa => yt_rsc_0_15_comp_qa,
      qb => yt_rsc_0_15_comp_qb,
      wea => yt_rsc_0_15_wea
    );
  yt_rsc_0_15_comp_adra <= yt_rsc_0_15_adra;
  yt_rsc_0_15_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_15_comp_da <= yt_rsc_0_15_da;
  yt_rsc_0_15_qa <= yt_rsc_0_15_comp_qa;
  yt_rsc_0_15_unc_1 <= yt_rsc_0_15_comp_qb;

  yt_rsc_0_16_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_16_comp_adra,
      adrb => yt_rsc_0_16_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_16_clken,
      da => yt_rsc_0_16_comp_da,
      qa => yt_rsc_0_16_comp_qa,
      qb => yt_rsc_0_16_comp_qb,
      wea => yt_rsc_0_16_wea
    );
  yt_rsc_0_16_comp_adra <= yt_rsc_0_16_adra;
  yt_rsc_0_16_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_16_comp_da <= yt_rsc_0_16_da;
  yt_rsc_0_16_qa <= yt_rsc_0_16_comp_qa;
  yt_rsc_0_16_unc_1 <= yt_rsc_0_16_comp_qb;

  yt_rsc_0_17_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_17_comp_adra,
      adrb => yt_rsc_0_17_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_17_clken,
      da => yt_rsc_0_17_comp_da,
      qa => yt_rsc_0_17_comp_qa,
      qb => yt_rsc_0_17_comp_qb,
      wea => yt_rsc_0_17_wea
    );
  yt_rsc_0_17_comp_adra <= yt_rsc_0_17_adra;
  yt_rsc_0_17_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_17_comp_da <= yt_rsc_0_17_da;
  yt_rsc_0_17_qa <= yt_rsc_0_17_comp_qa;
  yt_rsc_0_17_unc_1 <= yt_rsc_0_17_comp_qb;

  yt_rsc_0_18_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_18_comp_adra,
      adrb => yt_rsc_0_18_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_18_clken,
      da => yt_rsc_0_18_comp_da,
      qa => yt_rsc_0_18_comp_qa,
      qb => yt_rsc_0_18_comp_qb,
      wea => yt_rsc_0_18_wea
    );
  yt_rsc_0_18_comp_adra <= yt_rsc_0_18_adra;
  yt_rsc_0_18_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_18_comp_da <= yt_rsc_0_18_da;
  yt_rsc_0_18_qa <= yt_rsc_0_18_comp_qa;
  yt_rsc_0_18_unc_1 <= yt_rsc_0_18_comp_qb;

  yt_rsc_0_19_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_19_comp_adra,
      adrb => yt_rsc_0_19_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_19_clken,
      da => yt_rsc_0_19_comp_da,
      qa => yt_rsc_0_19_comp_qa,
      qb => yt_rsc_0_19_comp_qb,
      wea => yt_rsc_0_19_wea
    );
  yt_rsc_0_19_comp_adra <= yt_rsc_0_19_adra;
  yt_rsc_0_19_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_19_comp_da <= yt_rsc_0_19_da;
  yt_rsc_0_19_qa <= yt_rsc_0_19_comp_qa;
  yt_rsc_0_19_unc_1 <= yt_rsc_0_19_comp_qb;

  yt_rsc_0_20_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_20_comp_adra,
      adrb => yt_rsc_0_20_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_20_clken,
      da => yt_rsc_0_20_comp_da,
      qa => yt_rsc_0_20_comp_qa,
      qb => yt_rsc_0_20_comp_qb,
      wea => yt_rsc_0_20_wea
    );
  yt_rsc_0_20_comp_adra <= yt_rsc_0_20_adra;
  yt_rsc_0_20_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_20_comp_da <= yt_rsc_0_20_da;
  yt_rsc_0_20_qa <= yt_rsc_0_20_comp_qa;
  yt_rsc_0_20_unc_1 <= yt_rsc_0_20_comp_qb;

  yt_rsc_0_21_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_21_comp_adra,
      adrb => yt_rsc_0_21_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_21_clken,
      da => yt_rsc_0_21_comp_da,
      qa => yt_rsc_0_21_comp_qa,
      qb => yt_rsc_0_21_comp_qb,
      wea => yt_rsc_0_21_wea
    );
  yt_rsc_0_21_comp_adra <= yt_rsc_0_21_adra;
  yt_rsc_0_21_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_21_comp_da <= yt_rsc_0_21_da;
  yt_rsc_0_21_qa <= yt_rsc_0_21_comp_qa;
  yt_rsc_0_21_unc_1 <= yt_rsc_0_21_comp_qb;

  yt_rsc_0_22_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_22_comp_adra,
      adrb => yt_rsc_0_22_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_22_clken,
      da => yt_rsc_0_22_comp_da,
      qa => yt_rsc_0_22_comp_qa,
      qb => yt_rsc_0_22_comp_qb,
      wea => yt_rsc_0_22_wea
    );
  yt_rsc_0_22_comp_adra <= yt_rsc_0_22_adra;
  yt_rsc_0_22_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_22_comp_da <= yt_rsc_0_22_da;
  yt_rsc_0_22_qa <= yt_rsc_0_22_comp_qa;
  yt_rsc_0_22_unc_1 <= yt_rsc_0_22_comp_qb;

  yt_rsc_0_23_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_23_comp_adra,
      adrb => yt_rsc_0_23_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_23_clken,
      da => yt_rsc_0_23_comp_da,
      qa => yt_rsc_0_23_comp_qa,
      qb => yt_rsc_0_23_comp_qb,
      wea => yt_rsc_0_23_wea
    );
  yt_rsc_0_23_comp_adra <= yt_rsc_0_23_adra;
  yt_rsc_0_23_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_23_comp_da <= yt_rsc_0_23_da;
  yt_rsc_0_23_qa <= yt_rsc_0_23_comp_qa;
  yt_rsc_0_23_unc_1 <= yt_rsc_0_23_comp_qb;

  yt_rsc_0_24_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_24_comp_adra,
      adrb => yt_rsc_0_24_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_24_clken,
      da => yt_rsc_0_24_comp_da,
      qa => yt_rsc_0_24_comp_qa,
      qb => yt_rsc_0_24_comp_qb,
      wea => yt_rsc_0_24_wea
    );
  yt_rsc_0_24_comp_adra <= yt_rsc_0_24_adra;
  yt_rsc_0_24_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_24_comp_da <= yt_rsc_0_24_da;
  yt_rsc_0_24_qa <= yt_rsc_0_24_comp_qa;
  yt_rsc_0_24_unc_1 <= yt_rsc_0_24_comp_qb;

  yt_rsc_0_25_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_25_comp_adra,
      adrb => yt_rsc_0_25_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_25_clken,
      da => yt_rsc_0_25_comp_da,
      qa => yt_rsc_0_25_comp_qa,
      qb => yt_rsc_0_25_comp_qb,
      wea => yt_rsc_0_25_wea
    );
  yt_rsc_0_25_comp_adra <= yt_rsc_0_25_adra;
  yt_rsc_0_25_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_25_comp_da <= yt_rsc_0_25_da;
  yt_rsc_0_25_qa <= yt_rsc_0_25_comp_qa;
  yt_rsc_0_25_unc_1 <= yt_rsc_0_25_comp_qb;

  yt_rsc_0_26_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_26_comp_adra,
      adrb => yt_rsc_0_26_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_26_clken,
      da => yt_rsc_0_26_comp_da,
      qa => yt_rsc_0_26_comp_qa,
      qb => yt_rsc_0_26_comp_qb,
      wea => yt_rsc_0_26_wea
    );
  yt_rsc_0_26_comp_adra <= yt_rsc_0_26_adra;
  yt_rsc_0_26_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_26_comp_da <= yt_rsc_0_26_da;
  yt_rsc_0_26_qa <= yt_rsc_0_26_comp_qa;
  yt_rsc_0_26_unc_1 <= yt_rsc_0_26_comp_qb;

  yt_rsc_0_27_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_27_comp_adra,
      adrb => yt_rsc_0_27_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_27_clken,
      da => yt_rsc_0_27_comp_da,
      qa => yt_rsc_0_27_comp_qa,
      qb => yt_rsc_0_27_comp_qb,
      wea => yt_rsc_0_27_wea
    );
  yt_rsc_0_27_comp_adra <= yt_rsc_0_27_adra;
  yt_rsc_0_27_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_27_comp_da <= yt_rsc_0_27_da;
  yt_rsc_0_27_qa <= yt_rsc_0_27_comp_qa;
  yt_rsc_0_27_unc_1 <= yt_rsc_0_27_comp_qb;

  yt_rsc_0_28_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_28_comp_adra,
      adrb => yt_rsc_0_28_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_28_clken,
      da => yt_rsc_0_28_comp_da,
      qa => yt_rsc_0_28_comp_qa,
      qb => yt_rsc_0_28_comp_qb,
      wea => yt_rsc_0_28_wea
    );
  yt_rsc_0_28_comp_adra <= yt_rsc_0_28_adra;
  yt_rsc_0_28_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_28_comp_da <= yt_rsc_0_28_da;
  yt_rsc_0_28_qa <= yt_rsc_0_28_comp_qa;
  yt_rsc_0_28_unc_1 <= yt_rsc_0_28_comp_qb;

  yt_rsc_0_29_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_29_comp_adra,
      adrb => yt_rsc_0_29_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_29_clken,
      da => yt_rsc_0_29_comp_da,
      qa => yt_rsc_0_29_comp_qa,
      qb => yt_rsc_0_29_comp_qb,
      wea => yt_rsc_0_29_wea
    );
  yt_rsc_0_29_comp_adra <= yt_rsc_0_29_adra;
  yt_rsc_0_29_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_29_comp_da <= yt_rsc_0_29_da;
  yt_rsc_0_29_qa <= yt_rsc_0_29_comp_qa;
  yt_rsc_0_29_unc_1 <= yt_rsc_0_29_comp_qb;

  yt_rsc_0_30_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_30_comp_adra,
      adrb => yt_rsc_0_30_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_30_clken,
      da => yt_rsc_0_30_comp_da,
      qa => yt_rsc_0_30_comp_qa,
      qb => yt_rsc_0_30_comp_qb,
      wea => yt_rsc_0_30_wea
    );
  yt_rsc_0_30_comp_adra <= yt_rsc_0_30_adra;
  yt_rsc_0_30_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_30_comp_da <= yt_rsc_0_30_da;
  yt_rsc_0_30_qa <= yt_rsc_0_30_comp_qa;
  yt_rsc_0_30_unc_1 <= yt_rsc_0_30_comp_qb;

  yt_rsc_0_31_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_0_31_comp_adra,
      adrb => yt_rsc_0_31_comp_adrb,
      clk => clk,
      clken => yt_rsc_0_31_clken,
      da => yt_rsc_0_31_comp_da,
      qa => yt_rsc_0_31_comp_qa,
      qb => yt_rsc_0_31_comp_qb,
      wea => yt_rsc_0_31_wea
    );
  yt_rsc_0_31_comp_adra <= yt_rsc_0_31_adra;
  yt_rsc_0_31_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_0_31_comp_da <= yt_rsc_0_31_da;
  yt_rsc_0_31_qa <= yt_rsc_0_31_comp_qa;
  yt_rsc_0_31_unc_1 <= yt_rsc_0_31_comp_qb;

  yt_rsc_1_0_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_0_comp_adra,
      adrb => yt_rsc_1_0_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_0_clken,
      da => yt_rsc_1_0_comp_da,
      qa => yt_rsc_1_0_comp_qa,
      qb => yt_rsc_1_0_comp_qb,
      wea => yt_rsc_1_0_wea
    );
  yt_rsc_1_0_comp_adra <= yt_rsc_1_0_adra;
  yt_rsc_1_0_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_0_comp_da <= yt_rsc_1_0_da;
  yt_rsc_1_0_qa <= yt_rsc_1_0_comp_qa;
  yt_rsc_1_0_unc_1 <= yt_rsc_1_0_comp_qb;

  yt_rsc_1_1_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_1_comp_adra,
      adrb => yt_rsc_1_1_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_1_clken,
      da => yt_rsc_1_1_comp_da,
      qa => yt_rsc_1_1_comp_qa,
      qb => yt_rsc_1_1_comp_qb,
      wea => yt_rsc_1_1_wea
    );
  yt_rsc_1_1_comp_adra <= yt_rsc_1_1_adra;
  yt_rsc_1_1_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_1_comp_da <= yt_rsc_1_1_da;
  yt_rsc_1_1_qa <= yt_rsc_1_1_comp_qa;
  yt_rsc_1_1_unc_1 <= yt_rsc_1_1_comp_qb;

  yt_rsc_1_2_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_2_comp_adra,
      adrb => yt_rsc_1_2_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_2_clken,
      da => yt_rsc_1_2_comp_da,
      qa => yt_rsc_1_2_comp_qa,
      qb => yt_rsc_1_2_comp_qb,
      wea => yt_rsc_1_2_wea
    );
  yt_rsc_1_2_comp_adra <= yt_rsc_1_2_adra;
  yt_rsc_1_2_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_2_comp_da <= yt_rsc_1_2_da;
  yt_rsc_1_2_qa <= yt_rsc_1_2_comp_qa;
  yt_rsc_1_2_unc_1 <= yt_rsc_1_2_comp_qb;

  yt_rsc_1_3_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_3_comp_adra,
      adrb => yt_rsc_1_3_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_3_clken,
      da => yt_rsc_1_3_comp_da,
      qa => yt_rsc_1_3_comp_qa,
      qb => yt_rsc_1_3_comp_qb,
      wea => yt_rsc_1_3_wea
    );
  yt_rsc_1_3_comp_adra <= yt_rsc_1_3_adra;
  yt_rsc_1_3_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_3_comp_da <= yt_rsc_1_3_da;
  yt_rsc_1_3_qa <= yt_rsc_1_3_comp_qa;
  yt_rsc_1_3_unc_1 <= yt_rsc_1_3_comp_qb;

  yt_rsc_1_4_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_4_comp_adra,
      adrb => yt_rsc_1_4_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_4_clken,
      da => yt_rsc_1_4_comp_da,
      qa => yt_rsc_1_4_comp_qa,
      qb => yt_rsc_1_4_comp_qb,
      wea => yt_rsc_1_4_wea
    );
  yt_rsc_1_4_comp_adra <= yt_rsc_1_4_adra;
  yt_rsc_1_4_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_4_comp_da <= yt_rsc_1_4_da;
  yt_rsc_1_4_qa <= yt_rsc_1_4_comp_qa;
  yt_rsc_1_4_unc_1 <= yt_rsc_1_4_comp_qb;

  yt_rsc_1_5_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_5_comp_adra,
      adrb => yt_rsc_1_5_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_5_clken,
      da => yt_rsc_1_5_comp_da,
      qa => yt_rsc_1_5_comp_qa,
      qb => yt_rsc_1_5_comp_qb,
      wea => yt_rsc_1_5_wea
    );
  yt_rsc_1_5_comp_adra <= yt_rsc_1_5_adra;
  yt_rsc_1_5_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_5_comp_da <= yt_rsc_1_5_da;
  yt_rsc_1_5_qa <= yt_rsc_1_5_comp_qa;
  yt_rsc_1_5_unc_1 <= yt_rsc_1_5_comp_qb;

  yt_rsc_1_6_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_6_comp_adra,
      adrb => yt_rsc_1_6_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_6_clken,
      da => yt_rsc_1_6_comp_da,
      qa => yt_rsc_1_6_comp_qa,
      qb => yt_rsc_1_6_comp_qb,
      wea => yt_rsc_1_6_wea
    );
  yt_rsc_1_6_comp_adra <= yt_rsc_1_6_adra;
  yt_rsc_1_6_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_6_comp_da <= yt_rsc_1_6_da;
  yt_rsc_1_6_qa <= yt_rsc_1_6_comp_qa;
  yt_rsc_1_6_unc_1 <= yt_rsc_1_6_comp_qb;

  yt_rsc_1_7_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_7_comp_adra,
      adrb => yt_rsc_1_7_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_7_clken,
      da => yt_rsc_1_7_comp_da,
      qa => yt_rsc_1_7_comp_qa,
      qb => yt_rsc_1_7_comp_qb,
      wea => yt_rsc_1_7_wea
    );
  yt_rsc_1_7_comp_adra <= yt_rsc_1_7_adra;
  yt_rsc_1_7_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_7_comp_da <= yt_rsc_1_7_da;
  yt_rsc_1_7_qa <= yt_rsc_1_7_comp_qa;
  yt_rsc_1_7_unc_1 <= yt_rsc_1_7_comp_qb;

  yt_rsc_1_8_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_8_comp_adra,
      adrb => yt_rsc_1_8_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_8_clken,
      da => yt_rsc_1_8_comp_da,
      qa => yt_rsc_1_8_comp_qa,
      qb => yt_rsc_1_8_comp_qb,
      wea => yt_rsc_1_8_wea
    );
  yt_rsc_1_8_comp_adra <= yt_rsc_1_8_adra;
  yt_rsc_1_8_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_8_comp_da <= yt_rsc_1_8_da;
  yt_rsc_1_8_qa <= yt_rsc_1_8_comp_qa;
  yt_rsc_1_8_unc_1 <= yt_rsc_1_8_comp_qb;

  yt_rsc_1_9_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_9_comp_adra,
      adrb => yt_rsc_1_9_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_9_clken,
      da => yt_rsc_1_9_comp_da,
      qa => yt_rsc_1_9_comp_qa,
      qb => yt_rsc_1_9_comp_qb,
      wea => yt_rsc_1_9_wea
    );
  yt_rsc_1_9_comp_adra <= yt_rsc_1_9_adra;
  yt_rsc_1_9_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_9_comp_da <= yt_rsc_1_9_da;
  yt_rsc_1_9_qa <= yt_rsc_1_9_comp_qa;
  yt_rsc_1_9_unc_1 <= yt_rsc_1_9_comp_qb;

  yt_rsc_1_10_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_10_comp_adra,
      adrb => yt_rsc_1_10_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_10_clken,
      da => yt_rsc_1_10_comp_da,
      qa => yt_rsc_1_10_comp_qa,
      qb => yt_rsc_1_10_comp_qb,
      wea => yt_rsc_1_10_wea
    );
  yt_rsc_1_10_comp_adra <= yt_rsc_1_10_adra;
  yt_rsc_1_10_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_10_comp_da <= yt_rsc_1_10_da;
  yt_rsc_1_10_qa <= yt_rsc_1_10_comp_qa;
  yt_rsc_1_10_unc_1 <= yt_rsc_1_10_comp_qb;

  yt_rsc_1_11_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_11_comp_adra,
      adrb => yt_rsc_1_11_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_11_clken,
      da => yt_rsc_1_11_comp_da,
      qa => yt_rsc_1_11_comp_qa,
      qb => yt_rsc_1_11_comp_qb,
      wea => yt_rsc_1_11_wea
    );
  yt_rsc_1_11_comp_adra <= yt_rsc_1_11_adra;
  yt_rsc_1_11_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_11_comp_da <= yt_rsc_1_11_da;
  yt_rsc_1_11_qa <= yt_rsc_1_11_comp_qa;
  yt_rsc_1_11_unc_1 <= yt_rsc_1_11_comp_qb;

  yt_rsc_1_12_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_12_comp_adra,
      adrb => yt_rsc_1_12_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_12_clken,
      da => yt_rsc_1_12_comp_da,
      qa => yt_rsc_1_12_comp_qa,
      qb => yt_rsc_1_12_comp_qb,
      wea => yt_rsc_1_12_wea
    );
  yt_rsc_1_12_comp_adra <= yt_rsc_1_12_adra;
  yt_rsc_1_12_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_12_comp_da <= yt_rsc_1_12_da;
  yt_rsc_1_12_qa <= yt_rsc_1_12_comp_qa;
  yt_rsc_1_12_unc_1 <= yt_rsc_1_12_comp_qb;

  yt_rsc_1_13_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_13_comp_adra,
      adrb => yt_rsc_1_13_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_13_clken,
      da => yt_rsc_1_13_comp_da,
      qa => yt_rsc_1_13_comp_qa,
      qb => yt_rsc_1_13_comp_qb,
      wea => yt_rsc_1_13_wea
    );
  yt_rsc_1_13_comp_adra <= yt_rsc_1_13_adra;
  yt_rsc_1_13_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_13_comp_da <= yt_rsc_1_13_da;
  yt_rsc_1_13_qa <= yt_rsc_1_13_comp_qa;
  yt_rsc_1_13_unc_1 <= yt_rsc_1_13_comp_qb;

  yt_rsc_1_14_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_14_comp_adra,
      adrb => yt_rsc_1_14_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_14_clken,
      da => yt_rsc_1_14_comp_da,
      qa => yt_rsc_1_14_comp_qa,
      qb => yt_rsc_1_14_comp_qb,
      wea => yt_rsc_1_14_wea
    );
  yt_rsc_1_14_comp_adra <= yt_rsc_1_14_adra;
  yt_rsc_1_14_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_14_comp_da <= yt_rsc_1_14_da;
  yt_rsc_1_14_qa <= yt_rsc_1_14_comp_qa;
  yt_rsc_1_14_unc_1 <= yt_rsc_1_14_comp_qb;

  yt_rsc_1_15_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_15_comp_adra,
      adrb => yt_rsc_1_15_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_15_clken,
      da => yt_rsc_1_15_comp_da,
      qa => yt_rsc_1_15_comp_qa,
      qb => yt_rsc_1_15_comp_qb,
      wea => yt_rsc_1_15_wea
    );
  yt_rsc_1_15_comp_adra <= yt_rsc_1_15_adra;
  yt_rsc_1_15_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_15_comp_da <= yt_rsc_1_15_da;
  yt_rsc_1_15_qa <= yt_rsc_1_15_comp_qa;
  yt_rsc_1_15_unc_1 <= yt_rsc_1_15_comp_qb;

  yt_rsc_1_16_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_16_comp_adra,
      adrb => yt_rsc_1_16_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_16_clken,
      da => yt_rsc_1_16_comp_da,
      qa => yt_rsc_1_16_comp_qa,
      qb => yt_rsc_1_16_comp_qb,
      wea => yt_rsc_1_16_wea
    );
  yt_rsc_1_16_comp_adra <= yt_rsc_1_16_adra;
  yt_rsc_1_16_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_16_comp_da <= yt_rsc_1_16_da;
  yt_rsc_1_16_qa <= yt_rsc_1_16_comp_qa;
  yt_rsc_1_16_unc_1 <= yt_rsc_1_16_comp_qb;

  yt_rsc_1_17_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_17_comp_adra,
      adrb => yt_rsc_1_17_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_17_clken,
      da => yt_rsc_1_17_comp_da,
      qa => yt_rsc_1_17_comp_qa,
      qb => yt_rsc_1_17_comp_qb,
      wea => yt_rsc_1_17_wea
    );
  yt_rsc_1_17_comp_adra <= yt_rsc_1_17_adra;
  yt_rsc_1_17_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_17_comp_da <= yt_rsc_1_17_da;
  yt_rsc_1_17_qa <= yt_rsc_1_17_comp_qa;
  yt_rsc_1_17_unc_1 <= yt_rsc_1_17_comp_qb;

  yt_rsc_1_18_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_18_comp_adra,
      adrb => yt_rsc_1_18_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_18_clken,
      da => yt_rsc_1_18_comp_da,
      qa => yt_rsc_1_18_comp_qa,
      qb => yt_rsc_1_18_comp_qb,
      wea => yt_rsc_1_18_wea
    );
  yt_rsc_1_18_comp_adra <= yt_rsc_1_18_adra;
  yt_rsc_1_18_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_18_comp_da <= yt_rsc_1_18_da;
  yt_rsc_1_18_qa <= yt_rsc_1_18_comp_qa;
  yt_rsc_1_18_unc_1 <= yt_rsc_1_18_comp_qb;

  yt_rsc_1_19_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_19_comp_adra,
      adrb => yt_rsc_1_19_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_19_clken,
      da => yt_rsc_1_19_comp_da,
      qa => yt_rsc_1_19_comp_qa,
      qb => yt_rsc_1_19_comp_qb,
      wea => yt_rsc_1_19_wea
    );
  yt_rsc_1_19_comp_adra <= yt_rsc_1_19_adra;
  yt_rsc_1_19_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_19_comp_da <= yt_rsc_1_19_da;
  yt_rsc_1_19_qa <= yt_rsc_1_19_comp_qa;
  yt_rsc_1_19_unc_1 <= yt_rsc_1_19_comp_qb;

  yt_rsc_1_20_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_20_comp_adra,
      adrb => yt_rsc_1_20_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_20_clken,
      da => yt_rsc_1_20_comp_da,
      qa => yt_rsc_1_20_comp_qa,
      qb => yt_rsc_1_20_comp_qb,
      wea => yt_rsc_1_20_wea
    );
  yt_rsc_1_20_comp_adra <= yt_rsc_1_20_adra;
  yt_rsc_1_20_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_20_comp_da <= yt_rsc_1_20_da;
  yt_rsc_1_20_qa <= yt_rsc_1_20_comp_qa;
  yt_rsc_1_20_unc_1 <= yt_rsc_1_20_comp_qb;

  yt_rsc_1_21_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_21_comp_adra,
      adrb => yt_rsc_1_21_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_21_clken,
      da => yt_rsc_1_21_comp_da,
      qa => yt_rsc_1_21_comp_qa,
      qb => yt_rsc_1_21_comp_qb,
      wea => yt_rsc_1_21_wea
    );
  yt_rsc_1_21_comp_adra <= yt_rsc_1_21_adra;
  yt_rsc_1_21_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_21_comp_da <= yt_rsc_1_21_da;
  yt_rsc_1_21_qa <= yt_rsc_1_21_comp_qa;
  yt_rsc_1_21_unc_1 <= yt_rsc_1_21_comp_qb;

  yt_rsc_1_22_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_22_comp_adra,
      adrb => yt_rsc_1_22_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_22_clken,
      da => yt_rsc_1_22_comp_da,
      qa => yt_rsc_1_22_comp_qa,
      qb => yt_rsc_1_22_comp_qb,
      wea => yt_rsc_1_22_wea
    );
  yt_rsc_1_22_comp_adra <= yt_rsc_1_22_adra;
  yt_rsc_1_22_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_22_comp_da <= yt_rsc_1_22_da;
  yt_rsc_1_22_qa <= yt_rsc_1_22_comp_qa;
  yt_rsc_1_22_unc_1 <= yt_rsc_1_22_comp_qb;

  yt_rsc_1_23_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_23_comp_adra,
      adrb => yt_rsc_1_23_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_23_clken,
      da => yt_rsc_1_23_comp_da,
      qa => yt_rsc_1_23_comp_qa,
      qb => yt_rsc_1_23_comp_qb,
      wea => yt_rsc_1_23_wea
    );
  yt_rsc_1_23_comp_adra <= yt_rsc_1_23_adra;
  yt_rsc_1_23_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_23_comp_da <= yt_rsc_1_23_da;
  yt_rsc_1_23_qa <= yt_rsc_1_23_comp_qa;
  yt_rsc_1_23_unc_1 <= yt_rsc_1_23_comp_qb;

  yt_rsc_1_24_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_24_comp_adra,
      adrb => yt_rsc_1_24_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_24_clken,
      da => yt_rsc_1_24_comp_da,
      qa => yt_rsc_1_24_comp_qa,
      qb => yt_rsc_1_24_comp_qb,
      wea => yt_rsc_1_24_wea
    );
  yt_rsc_1_24_comp_adra <= yt_rsc_1_24_adra;
  yt_rsc_1_24_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_24_comp_da <= yt_rsc_1_24_da;
  yt_rsc_1_24_qa <= yt_rsc_1_24_comp_qa;
  yt_rsc_1_24_unc_1 <= yt_rsc_1_24_comp_qb;

  yt_rsc_1_25_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_25_comp_adra,
      adrb => yt_rsc_1_25_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_25_clken,
      da => yt_rsc_1_25_comp_da,
      qa => yt_rsc_1_25_comp_qa,
      qb => yt_rsc_1_25_comp_qb,
      wea => yt_rsc_1_25_wea
    );
  yt_rsc_1_25_comp_adra <= yt_rsc_1_25_adra;
  yt_rsc_1_25_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_25_comp_da <= yt_rsc_1_25_da;
  yt_rsc_1_25_qa <= yt_rsc_1_25_comp_qa;
  yt_rsc_1_25_unc_1 <= yt_rsc_1_25_comp_qb;

  yt_rsc_1_26_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_26_comp_adra,
      adrb => yt_rsc_1_26_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_26_clken,
      da => yt_rsc_1_26_comp_da,
      qa => yt_rsc_1_26_comp_qa,
      qb => yt_rsc_1_26_comp_qb,
      wea => yt_rsc_1_26_wea
    );
  yt_rsc_1_26_comp_adra <= yt_rsc_1_26_adra;
  yt_rsc_1_26_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_26_comp_da <= yt_rsc_1_26_da;
  yt_rsc_1_26_qa <= yt_rsc_1_26_comp_qa;
  yt_rsc_1_26_unc_1 <= yt_rsc_1_26_comp_qb;

  yt_rsc_1_27_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_27_comp_adra,
      adrb => yt_rsc_1_27_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_27_clken,
      da => yt_rsc_1_27_comp_da,
      qa => yt_rsc_1_27_comp_qa,
      qb => yt_rsc_1_27_comp_qb,
      wea => yt_rsc_1_27_wea
    );
  yt_rsc_1_27_comp_adra <= yt_rsc_1_27_adra;
  yt_rsc_1_27_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_27_comp_da <= yt_rsc_1_27_da;
  yt_rsc_1_27_qa <= yt_rsc_1_27_comp_qa;
  yt_rsc_1_27_unc_1 <= yt_rsc_1_27_comp_qb;

  yt_rsc_1_28_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_28_comp_adra,
      adrb => yt_rsc_1_28_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_28_clken,
      da => yt_rsc_1_28_comp_da,
      qa => yt_rsc_1_28_comp_qa,
      qb => yt_rsc_1_28_comp_qb,
      wea => yt_rsc_1_28_wea
    );
  yt_rsc_1_28_comp_adra <= yt_rsc_1_28_adra;
  yt_rsc_1_28_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_28_comp_da <= yt_rsc_1_28_da;
  yt_rsc_1_28_qa <= yt_rsc_1_28_comp_qa;
  yt_rsc_1_28_unc_1 <= yt_rsc_1_28_comp_qb;

  yt_rsc_1_29_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_29_comp_adra,
      adrb => yt_rsc_1_29_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_29_clken,
      da => yt_rsc_1_29_comp_da,
      qa => yt_rsc_1_29_comp_qa,
      qb => yt_rsc_1_29_comp_qb,
      wea => yt_rsc_1_29_wea
    );
  yt_rsc_1_29_comp_adra <= yt_rsc_1_29_adra;
  yt_rsc_1_29_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_29_comp_da <= yt_rsc_1_29_da;
  yt_rsc_1_29_qa <= yt_rsc_1_29_comp_qa;
  yt_rsc_1_29_unc_1 <= yt_rsc_1_29_comp_qb;

  yt_rsc_1_30_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_30_comp_adra,
      adrb => yt_rsc_1_30_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_30_clken,
      da => yt_rsc_1_30_comp_da,
      qa => yt_rsc_1_30_comp_qa,
      qb => yt_rsc_1_30_comp_qb,
      wea => yt_rsc_1_30_wea
    );
  yt_rsc_1_30_comp_adra <= yt_rsc_1_30_adra;
  yt_rsc_1_30_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_30_comp_da <= yt_rsc_1_30_da;
  yt_rsc_1_30_qa <= yt_rsc_1_30_comp_qa;
  yt_rsc_1_30_unc_1 <= yt_rsc_1_30_comp_qb;

  yt_rsc_1_31_comp : work.block_2r1w_rbw_pkg.BLOCK_2R1W_RBW
    GENERIC MAP(
      addr_width => 4,
      data_width => 32,
      depth => 16,
      latency => 1
      )
    PORT MAP(
      adra => yt_rsc_1_31_comp_adra,
      adrb => yt_rsc_1_31_comp_adrb,
      clk => clk,
      clken => yt_rsc_1_31_clken,
      da => yt_rsc_1_31_comp_da,
      qa => yt_rsc_1_31_comp_qa,
      qb => yt_rsc_1_31_comp_qb,
      wea => yt_rsc_1_31_wea
    );
  yt_rsc_1_31_comp_adra <= yt_rsc_1_31_adra;
  yt_rsc_1_31_comp_adrb <= STD_LOGIC_VECTOR'( "0000");
  yt_rsc_1_31_comp_da <= yt_rsc_1_31_da;
  yt_rsc_1_31_qa <= yt_rsc_1_31_comp_qa;
  yt_rsc_1_31_unc_1 <= yt_rsc_1_31_comp_qb;

  yt_rsc_0_0_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_7_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_0_clken,
      qa => yt_rsc_0_0_i_qa,
      wea => yt_rsc_0_0_wea,
      da => yt_rsc_0_0_i_da,
      adra => yt_rsc_0_0_i_adra,
      adra_d => yt_rsc_0_0_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_0_i_da_d,
      qa_d => yt_rsc_0_0_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_0_i_qa <= yt_rsc_0_0_qa;
  yt_rsc_0_0_da <= yt_rsc_0_0_i_da;
  yt_rsc_0_0_adra <= yt_rsc_0_0_i_adra;
  yt_rsc_0_0_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_0_i_da_d <= yt_rsc_0_0_i_da_d_iff;
  yt_rsc_0_0_i_qa_d <= yt_rsc_0_0_i_qa_d_1;

  yt_rsc_0_1_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_8_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_1_clken,
      qa => yt_rsc_0_1_i_qa,
      wea => yt_rsc_0_1_wea,
      da => yt_rsc_0_1_i_da,
      adra => yt_rsc_0_1_i_adra,
      adra_d => yt_rsc_0_1_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_1_i_da_d,
      qa_d => yt_rsc_0_1_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_1_i_qa <= yt_rsc_0_1_qa;
  yt_rsc_0_1_da <= yt_rsc_0_1_i_da;
  yt_rsc_0_1_adra <= yt_rsc_0_1_i_adra;
  yt_rsc_0_1_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_1_i_da_d <= yt_rsc_0_1_i_da_d_iff;
  yt_rsc_0_1_i_qa_d <= yt_rsc_0_1_i_qa_d_1;

  yt_rsc_0_2_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_9_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_2_clken,
      qa => yt_rsc_0_2_i_qa,
      wea => yt_rsc_0_2_wea,
      da => yt_rsc_0_2_i_da,
      adra => yt_rsc_0_2_i_adra,
      adra_d => yt_rsc_0_2_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_2_i_da_d,
      qa_d => yt_rsc_0_2_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_2_i_qa <= yt_rsc_0_2_qa;
  yt_rsc_0_2_da <= yt_rsc_0_2_i_da;
  yt_rsc_0_2_adra <= yt_rsc_0_2_i_adra;
  yt_rsc_0_2_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_2_i_da_d <= yt_rsc_0_2_i_da_d_iff;
  yt_rsc_0_2_i_qa_d <= yt_rsc_0_2_i_qa_d_1;

  yt_rsc_0_3_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_10_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_3_clken,
      qa => yt_rsc_0_3_i_qa,
      wea => yt_rsc_0_3_wea,
      da => yt_rsc_0_3_i_da,
      adra => yt_rsc_0_3_i_adra,
      adra_d => yt_rsc_0_3_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_3_i_da_d,
      qa_d => yt_rsc_0_3_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_3_i_qa <= yt_rsc_0_3_qa;
  yt_rsc_0_3_da <= yt_rsc_0_3_i_da;
  yt_rsc_0_3_adra <= yt_rsc_0_3_i_adra;
  yt_rsc_0_3_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_3_i_da_d <= yt_rsc_0_3_i_da_d_iff;
  yt_rsc_0_3_i_qa_d <= yt_rsc_0_3_i_qa_d_1;

  yt_rsc_0_4_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_11_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_4_clken,
      qa => yt_rsc_0_4_i_qa,
      wea => yt_rsc_0_4_wea,
      da => yt_rsc_0_4_i_da,
      adra => yt_rsc_0_4_i_adra,
      adra_d => yt_rsc_0_4_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_4_i_da_d,
      qa_d => yt_rsc_0_4_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_4_i_qa <= yt_rsc_0_4_qa;
  yt_rsc_0_4_da <= yt_rsc_0_4_i_da;
  yt_rsc_0_4_adra <= yt_rsc_0_4_i_adra;
  yt_rsc_0_4_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_4_i_da_d <= yt_rsc_0_4_i_da_d_iff;
  yt_rsc_0_4_i_qa_d <= yt_rsc_0_4_i_qa_d_1;

  yt_rsc_0_5_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_12_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_5_clken,
      qa => yt_rsc_0_5_i_qa,
      wea => yt_rsc_0_5_wea,
      da => yt_rsc_0_5_i_da,
      adra => yt_rsc_0_5_i_adra,
      adra_d => yt_rsc_0_5_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_5_i_da_d,
      qa_d => yt_rsc_0_5_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_5_i_qa <= yt_rsc_0_5_qa;
  yt_rsc_0_5_da <= yt_rsc_0_5_i_da;
  yt_rsc_0_5_adra <= yt_rsc_0_5_i_adra;
  yt_rsc_0_5_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_5_i_da_d <= yt_rsc_0_5_i_da_d_iff;
  yt_rsc_0_5_i_qa_d <= yt_rsc_0_5_i_qa_d_1;

  yt_rsc_0_6_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_13_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_6_clken,
      qa => yt_rsc_0_6_i_qa,
      wea => yt_rsc_0_6_wea,
      da => yt_rsc_0_6_i_da,
      adra => yt_rsc_0_6_i_adra,
      adra_d => yt_rsc_0_6_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_6_i_da_d,
      qa_d => yt_rsc_0_6_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_6_i_qa <= yt_rsc_0_6_qa;
  yt_rsc_0_6_da <= yt_rsc_0_6_i_da;
  yt_rsc_0_6_adra <= yt_rsc_0_6_i_adra;
  yt_rsc_0_6_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_6_i_da_d <= yt_rsc_0_6_i_da_d_iff;
  yt_rsc_0_6_i_qa_d <= yt_rsc_0_6_i_qa_d_1;

  yt_rsc_0_7_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_14_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_7_clken,
      qa => yt_rsc_0_7_i_qa,
      wea => yt_rsc_0_7_wea,
      da => yt_rsc_0_7_i_da,
      adra => yt_rsc_0_7_i_adra,
      adra_d => yt_rsc_0_7_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_7_i_da_d,
      qa_d => yt_rsc_0_7_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_7_i_qa <= yt_rsc_0_7_qa;
  yt_rsc_0_7_da <= yt_rsc_0_7_i_da;
  yt_rsc_0_7_adra <= yt_rsc_0_7_i_adra;
  yt_rsc_0_7_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_7_i_da_d <= yt_rsc_0_7_i_da_d_iff;
  yt_rsc_0_7_i_qa_d <= yt_rsc_0_7_i_qa_d_1;

  yt_rsc_0_8_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_15_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_8_clken,
      qa => yt_rsc_0_8_i_qa,
      wea => yt_rsc_0_8_wea,
      da => yt_rsc_0_8_i_da,
      adra => yt_rsc_0_8_i_adra,
      adra_d => yt_rsc_0_8_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_8_i_da_d,
      qa_d => yt_rsc_0_8_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_8_i_qa <= yt_rsc_0_8_qa;
  yt_rsc_0_8_da <= yt_rsc_0_8_i_da;
  yt_rsc_0_8_adra <= yt_rsc_0_8_i_adra;
  yt_rsc_0_8_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_8_i_da_d <= yt_rsc_0_8_i_da_d_iff;
  yt_rsc_0_8_i_qa_d <= yt_rsc_0_8_i_qa_d_1;

  yt_rsc_0_9_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_16_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_9_clken,
      qa => yt_rsc_0_9_i_qa,
      wea => yt_rsc_0_9_wea,
      da => yt_rsc_0_9_i_da,
      adra => yt_rsc_0_9_i_adra,
      adra_d => yt_rsc_0_9_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_9_i_da_d,
      qa_d => yt_rsc_0_9_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_9_i_qa <= yt_rsc_0_9_qa;
  yt_rsc_0_9_da <= yt_rsc_0_9_i_da;
  yt_rsc_0_9_adra <= yt_rsc_0_9_i_adra;
  yt_rsc_0_9_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_9_i_da_d <= yt_rsc_0_9_i_da_d_iff;
  yt_rsc_0_9_i_qa_d <= yt_rsc_0_9_i_qa_d_1;

  yt_rsc_0_10_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_17_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_10_clken,
      qa => yt_rsc_0_10_i_qa,
      wea => yt_rsc_0_10_wea,
      da => yt_rsc_0_10_i_da,
      adra => yt_rsc_0_10_i_adra,
      adra_d => yt_rsc_0_10_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_10_i_da_d,
      qa_d => yt_rsc_0_10_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_10_i_qa <= yt_rsc_0_10_qa;
  yt_rsc_0_10_da <= yt_rsc_0_10_i_da;
  yt_rsc_0_10_adra <= yt_rsc_0_10_i_adra;
  yt_rsc_0_10_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_10_i_da_d <= yt_rsc_0_10_i_da_d_iff;
  yt_rsc_0_10_i_qa_d <= yt_rsc_0_10_i_qa_d_1;

  yt_rsc_0_11_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_18_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_11_clken,
      qa => yt_rsc_0_11_i_qa,
      wea => yt_rsc_0_11_wea,
      da => yt_rsc_0_11_i_da,
      adra => yt_rsc_0_11_i_adra,
      adra_d => yt_rsc_0_11_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_11_i_da_d,
      qa_d => yt_rsc_0_11_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_11_i_qa <= yt_rsc_0_11_qa;
  yt_rsc_0_11_da <= yt_rsc_0_11_i_da;
  yt_rsc_0_11_adra <= yt_rsc_0_11_i_adra;
  yt_rsc_0_11_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_11_i_da_d <= yt_rsc_0_11_i_da_d_iff;
  yt_rsc_0_11_i_qa_d <= yt_rsc_0_11_i_qa_d_1;

  yt_rsc_0_12_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_19_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_12_clken,
      qa => yt_rsc_0_12_i_qa,
      wea => yt_rsc_0_12_wea,
      da => yt_rsc_0_12_i_da,
      adra => yt_rsc_0_12_i_adra,
      adra_d => yt_rsc_0_12_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_12_i_da_d,
      qa_d => yt_rsc_0_12_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_12_i_qa <= yt_rsc_0_12_qa;
  yt_rsc_0_12_da <= yt_rsc_0_12_i_da;
  yt_rsc_0_12_adra <= yt_rsc_0_12_i_adra;
  yt_rsc_0_12_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_12_i_da_d <= yt_rsc_0_12_i_da_d_iff;
  yt_rsc_0_12_i_qa_d <= yt_rsc_0_12_i_qa_d_1;

  yt_rsc_0_13_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_20_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_13_clken,
      qa => yt_rsc_0_13_i_qa,
      wea => yt_rsc_0_13_wea,
      da => yt_rsc_0_13_i_da,
      adra => yt_rsc_0_13_i_adra,
      adra_d => yt_rsc_0_13_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_13_i_da_d,
      qa_d => yt_rsc_0_13_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_13_i_qa <= yt_rsc_0_13_qa;
  yt_rsc_0_13_da <= yt_rsc_0_13_i_da;
  yt_rsc_0_13_adra <= yt_rsc_0_13_i_adra;
  yt_rsc_0_13_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_13_i_da_d <= yt_rsc_0_13_i_da_d_iff;
  yt_rsc_0_13_i_qa_d <= yt_rsc_0_13_i_qa_d_1;

  yt_rsc_0_14_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_21_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_14_clken,
      qa => yt_rsc_0_14_i_qa,
      wea => yt_rsc_0_14_wea,
      da => yt_rsc_0_14_i_da,
      adra => yt_rsc_0_14_i_adra,
      adra_d => yt_rsc_0_14_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_14_i_da_d,
      qa_d => yt_rsc_0_14_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_14_i_qa <= yt_rsc_0_14_qa;
  yt_rsc_0_14_da <= yt_rsc_0_14_i_da;
  yt_rsc_0_14_adra <= yt_rsc_0_14_i_adra;
  yt_rsc_0_14_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_14_i_da_d <= yt_rsc_0_14_i_da_d_iff;
  yt_rsc_0_14_i_qa_d <= yt_rsc_0_14_i_qa_d_1;

  yt_rsc_0_15_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_22_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_15_clken,
      qa => yt_rsc_0_15_i_qa,
      wea => yt_rsc_0_15_wea,
      da => yt_rsc_0_15_i_da,
      adra => yt_rsc_0_15_i_adra,
      adra_d => yt_rsc_0_15_i_adra_d,
      clken_d => yt_rsc_0_0_i_clken_d,
      da_d => yt_rsc_0_15_i_da_d,
      qa_d => yt_rsc_0_15_i_qa_d_1,
      wea_d => yt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_0_i_wea_d_iff
    );
  yt_rsc_0_15_i_qa <= yt_rsc_0_15_qa;
  yt_rsc_0_15_da <= yt_rsc_0_15_i_da;
  yt_rsc_0_15_adra <= yt_rsc_0_15_i_adra;
  yt_rsc_0_15_i_adra_d <= yt_rsc_0_0_i_adra_d_iff;
  yt_rsc_0_15_i_da_d <= yt_rsc_0_15_i_da_d_iff;
  yt_rsc_0_15_i_qa_d <= yt_rsc_0_15_i_qa_d_1;

  yt_rsc_0_16_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_23_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_16_clken,
      qa => yt_rsc_0_16_i_qa,
      wea => yt_rsc_0_16_wea,
      da => yt_rsc_0_16_i_da,
      adra => yt_rsc_0_16_i_adra,
      adra_d => yt_rsc_0_16_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_16_i_da_d,
      qa_d => yt_rsc_0_16_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_16_i_qa <= yt_rsc_0_16_qa;
  yt_rsc_0_16_da <= yt_rsc_0_16_i_da;
  yt_rsc_0_16_adra <= yt_rsc_0_16_i_adra;
  yt_rsc_0_16_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_16_i_da_d <= yt_rsc_0_0_i_da_d_iff;
  yt_rsc_0_16_i_qa_d <= yt_rsc_0_16_i_qa_d_1;

  yt_rsc_0_17_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_24_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_17_clken,
      qa => yt_rsc_0_17_i_qa,
      wea => yt_rsc_0_17_wea,
      da => yt_rsc_0_17_i_da,
      adra => yt_rsc_0_17_i_adra,
      adra_d => yt_rsc_0_17_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_17_i_da_d,
      qa_d => yt_rsc_0_17_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_17_i_qa <= yt_rsc_0_17_qa;
  yt_rsc_0_17_da <= yt_rsc_0_17_i_da;
  yt_rsc_0_17_adra <= yt_rsc_0_17_i_adra;
  yt_rsc_0_17_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_17_i_da_d <= yt_rsc_0_1_i_da_d_iff;
  yt_rsc_0_17_i_qa_d <= yt_rsc_0_17_i_qa_d_1;

  yt_rsc_0_18_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_25_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_18_clken,
      qa => yt_rsc_0_18_i_qa,
      wea => yt_rsc_0_18_wea,
      da => yt_rsc_0_18_i_da,
      adra => yt_rsc_0_18_i_adra,
      adra_d => yt_rsc_0_18_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_18_i_da_d,
      qa_d => yt_rsc_0_18_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_18_i_qa <= yt_rsc_0_18_qa;
  yt_rsc_0_18_da <= yt_rsc_0_18_i_da;
  yt_rsc_0_18_adra <= yt_rsc_0_18_i_adra;
  yt_rsc_0_18_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_18_i_da_d <= yt_rsc_0_2_i_da_d_iff;
  yt_rsc_0_18_i_qa_d <= yt_rsc_0_18_i_qa_d_1;

  yt_rsc_0_19_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_26_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_19_clken,
      qa => yt_rsc_0_19_i_qa,
      wea => yt_rsc_0_19_wea,
      da => yt_rsc_0_19_i_da,
      adra => yt_rsc_0_19_i_adra,
      adra_d => yt_rsc_0_19_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_19_i_da_d,
      qa_d => yt_rsc_0_19_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_19_i_qa <= yt_rsc_0_19_qa;
  yt_rsc_0_19_da <= yt_rsc_0_19_i_da;
  yt_rsc_0_19_adra <= yt_rsc_0_19_i_adra;
  yt_rsc_0_19_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_19_i_da_d <= yt_rsc_0_3_i_da_d_iff;
  yt_rsc_0_19_i_qa_d <= yt_rsc_0_19_i_qa_d_1;

  yt_rsc_0_20_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_27_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_20_clken,
      qa => yt_rsc_0_20_i_qa,
      wea => yt_rsc_0_20_wea,
      da => yt_rsc_0_20_i_da,
      adra => yt_rsc_0_20_i_adra,
      adra_d => yt_rsc_0_20_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_20_i_da_d,
      qa_d => yt_rsc_0_20_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_20_i_qa <= yt_rsc_0_20_qa;
  yt_rsc_0_20_da <= yt_rsc_0_20_i_da;
  yt_rsc_0_20_adra <= yt_rsc_0_20_i_adra;
  yt_rsc_0_20_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_20_i_da_d <= yt_rsc_0_4_i_da_d_iff;
  yt_rsc_0_20_i_qa_d <= yt_rsc_0_20_i_qa_d_1;

  yt_rsc_0_21_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_28_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_21_clken,
      qa => yt_rsc_0_21_i_qa,
      wea => yt_rsc_0_21_wea,
      da => yt_rsc_0_21_i_da,
      adra => yt_rsc_0_21_i_adra,
      adra_d => yt_rsc_0_21_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_21_i_da_d,
      qa_d => yt_rsc_0_21_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_21_i_qa <= yt_rsc_0_21_qa;
  yt_rsc_0_21_da <= yt_rsc_0_21_i_da;
  yt_rsc_0_21_adra <= yt_rsc_0_21_i_adra;
  yt_rsc_0_21_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_21_i_da_d <= yt_rsc_0_5_i_da_d_iff;
  yt_rsc_0_21_i_qa_d <= yt_rsc_0_21_i_qa_d_1;

  yt_rsc_0_22_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_29_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_22_clken,
      qa => yt_rsc_0_22_i_qa,
      wea => yt_rsc_0_22_wea,
      da => yt_rsc_0_22_i_da,
      adra => yt_rsc_0_22_i_adra,
      adra_d => yt_rsc_0_22_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_22_i_da_d,
      qa_d => yt_rsc_0_22_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_22_i_qa <= yt_rsc_0_22_qa;
  yt_rsc_0_22_da <= yt_rsc_0_22_i_da;
  yt_rsc_0_22_adra <= yt_rsc_0_22_i_adra;
  yt_rsc_0_22_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_22_i_da_d <= yt_rsc_0_6_i_da_d_iff;
  yt_rsc_0_22_i_qa_d <= yt_rsc_0_22_i_qa_d_1;

  yt_rsc_0_23_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_30_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_23_clken,
      qa => yt_rsc_0_23_i_qa,
      wea => yt_rsc_0_23_wea,
      da => yt_rsc_0_23_i_da,
      adra => yt_rsc_0_23_i_adra,
      adra_d => yt_rsc_0_23_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_23_i_da_d,
      qa_d => yt_rsc_0_23_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_23_i_qa <= yt_rsc_0_23_qa;
  yt_rsc_0_23_da <= yt_rsc_0_23_i_da;
  yt_rsc_0_23_adra <= yt_rsc_0_23_i_adra;
  yt_rsc_0_23_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_23_i_da_d <= yt_rsc_0_7_i_da_d_iff;
  yt_rsc_0_23_i_qa_d <= yt_rsc_0_23_i_qa_d_1;

  yt_rsc_0_24_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_31_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_24_clken,
      qa => yt_rsc_0_24_i_qa,
      wea => yt_rsc_0_24_wea,
      da => yt_rsc_0_24_i_da,
      adra => yt_rsc_0_24_i_adra,
      adra_d => yt_rsc_0_24_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_24_i_da_d,
      qa_d => yt_rsc_0_24_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_24_i_qa <= yt_rsc_0_24_qa;
  yt_rsc_0_24_da <= yt_rsc_0_24_i_da;
  yt_rsc_0_24_adra <= yt_rsc_0_24_i_adra;
  yt_rsc_0_24_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_24_i_da_d <= yt_rsc_0_8_i_da_d_iff;
  yt_rsc_0_24_i_qa_d <= yt_rsc_0_24_i_qa_d_1;

  yt_rsc_0_25_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_32_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_25_clken,
      qa => yt_rsc_0_25_i_qa,
      wea => yt_rsc_0_25_wea,
      da => yt_rsc_0_25_i_da,
      adra => yt_rsc_0_25_i_adra,
      adra_d => yt_rsc_0_25_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_25_i_da_d,
      qa_d => yt_rsc_0_25_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_25_i_qa <= yt_rsc_0_25_qa;
  yt_rsc_0_25_da <= yt_rsc_0_25_i_da;
  yt_rsc_0_25_adra <= yt_rsc_0_25_i_adra;
  yt_rsc_0_25_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_25_i_da_d <= yt_rsc_0_9_i_da_d_iff;
  yt_rsc_0_25_i_qa_d <= yt_rsc_0_25_i_qa_d_1;

  yt_rsc_0_26_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_33_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_26_clken,
      qa => yt_rsc_0_26_i_qa,
      wea => yt_rsc_0_26_wea,
      da => yt_rsc_0_26_i_da,
      adra => yt_rsc_0_26_i_adra,
      adra_d => yt_rsc_0_26_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_26_i_da_d,
      qa_d => yt_rsc_0_26_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_26_i_qa <= yt_rsc_0_26_qa;
  yt_rsc_0_26_da <= yt_rsc_0_26_i_da;
  yt_rsc_0_26_adra <= yt_rsc_0_26_i_adra;
  yt_rsc_0_26_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_26_i_da_d <= yt_rsc_0_10_i_da_d_iff;
  yt_rsc_0_26_i_qa_d <= yt_rsc_0_26_i_qa_d_1;

  yt_rsc_0_27_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_34_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_27_clken,
      qa => yt_rsc_0_27_i_qa,
      wea => yt_rsc_0_27_wea,
      da => yt_rsc_0_27_i_da,
      adra => yt_rsc_0_27_i_adra,
      adra_d => yt_rsc_0_27_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_27_i_da_d,
      qa_d => yt_rsc_0_27_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_27_i_qa <= yt_rsc_0_27_qa;
  yt_rsc_0_27_da <= yt_rsc_0_27_i_da;
  yt_rsc_0_27_adra <= yt_rsc_0_27_i_adra;
  yt_rsc_0_27_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_27_i_da_d <= yt_rsc_0_11_i_da_d_iff;
  yt_rsc_0_27_i_qa_d <= yt_rsc_0_27_i_qa_d_1;

  yt_rsc_0_28_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_35_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_28_clken,
      qa => yt_rsc_0_28_i_qa,
      wea => yt_rsc_0_28_wea,
      da => yt_rsc_0_28_i_da,
      adra => yt_rsc_0_28_i_adra,
      adra_d => yt_rsc_0_28_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_28_i_da_d,
      qa_d => yt_rsc_0_28_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_28_i_qa <= yt_rsc_0_28_qa;
  yt_rsc_0_28_da <= yt_rsc_0_28_i_da;
  yt_rsc_0_28_adra <= yt_rsc_0_28_i_adra;
  yt_rsc_0_28_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_28_i_da_d <= yt_rsc_0_12_i_da_d_iff;
  yt_rsc_0_28_i_qa_d <= yt_rsc_0_28_i_qa_d_1;

  yt_rsc_0_29_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_36_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_29_clken,
      qa => yt_rsc_0_29_i_qa,
      wea => yt_rsc_0_29_wea,
      da => yt_rsc_0_29_i_da,
      adra => yt_rsc_0_29_i_adra,
      adra_d => yt_rsc_0_29_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_29_i_da_d,
      qa_d => yt_rsc_0_29_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_29_i_qa <= yt_rsc_0_29_qa;
  yt_rsc_0_29_da <= yt_rsc_0_29_i_da;
  yt_rsc_0_29_adra <= yt_rsc_0_29_i_adra;
  yt_rsc_0_29_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_29_i_da_d <= yt_rsc_0_13_i_da_d_iff;
  yt_rsc_0_29_i_qa_d <= yt_rsc_0_29_i_qa_d_1;

  yt_rsc_0_30_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_37_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_30_clken,
      qa => yt_rsc_0_30_i_qa,
      wea => yt_rsc_0_30_wea,
      da => yt_rsc_0_30_i_da,
      adra => yt_rsc_0_30_i_adra,
      adra_d => yt_rsc_0_30_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_30_i_da_d,
      qa_d => yt_rsc_0_30_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_30_i_qa <= yt_rsc_0_30_qa;
  yt_rsc_0_30_da <= yt_rsc_0_30_i_da;
  yt_rsc_0_30_adra <= yt_rsc_0_30_i_adra;
  yt_rsc_0_30_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_30_i_da_d <= yt_rsc_0_14_i_da_d_iff;
  yt_rsc_0_30_i_qa_d <= yt_rsc_0_30_i_qa_d_1;

  yt_rsc_0_31_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_38_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_0_31_clken,
      qa => yt_rsc_0_31_i_qa,
      wea => yt_rsc_0_31_wea,
      da => yt_rsc_0_31_i_da,
      adra => yt_rsc_0_31_i_adra,
      adra_d => yt_rsc_0_31_i_adra_d,
      clken_d => yt_rsc_0_16_i_clken_d,
      da_d => yt_rsc_0_31_i_da_d,
      qa_d => yt_rsc_0_31_i_qa_d_1,
      wea_d => yt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_0_16_i_wea_d_iff
    );
  yt_rsc_0_31_i_qa <= yt_rsc_0_31_qa;
  yt_rsc_0_31_da <= yt_rsc_0_31_i_da;
  yt_rsc_0_31_adra <= yt_rsc_0_31_i_adra;
  yt_rsc_0_31_i_adra_d <= yt_rsc_0_16_i_adra_d_iff;
  yt_rsc_0_31_i_da_d <= yt_rsc_0_15_i_da_d_iff;
  yt_rsc_0_31_i_qa_d <= yt_rsc_0_31_i_qa_d_1;

  yt_rsc_1_0_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_39_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_0_clken,
      qa => yt_rsc_1_0_i_qa,
      wea => yt_rsc_1_0_wea,
      da => yt_rsc_1_0_i_da,
      adra => yt_rsc_1_0_i_adra,
      adra_d => yt_rsc_1_0_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_0_i_da_d_1,
      qa_d => yt_rsc_1_0_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_0_i_qa <= yt_rsc_1_0_qa;
  yt_rsc_1_0_da <= yt_rsc_1_0_i_da;
  yt_rsc_1_0_adra <= yt_rsc_1_0_i_adra;
  yt_rsc_1_0_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_0_i_da_d_1 <= yt_rsc_1_0_i_da_d;
  yt_rsc_1_0_i_qa_d <= yt_rsc_1_0_i_qa_d_1;

  yt_rsc_1_1_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_40_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_1_clken,
      qa => yt_rsc_1_1_i_qa,
      wea => yt_rsc_1_1_wea,
      da => yt_rsc_1_1_i_da,
      adra => yt_rsc_1_1_i_adra,
      adra_d => yt_rsc_1_1_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_1_i_da_d_1,
      qa_d => yt_rsc_1_1_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_1_i_qa <= yt_rsc_1_1_qa;
  yt_rsc_1_1_da <= yt_rsc_1_1_i_da;
  yt_rsc_1_1_adra <= yt_rsc_1_1_i_adra;
  yt_rsc_1_1_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_1_i_da_d_1 <= yt_rsc_1_1_i_da_d;
  yt_rsc_1_1_i_qa_d <= yt_rsc_1_1_i_qa_d_1;

  yt_rsc_1_2_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_41_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_2_clken,
      qa => yt_rsc_1_2_i_qa,
      wea => yt_rsc_1_2_wea,
      da => yt_rsc_1_2_i_da,
      adra => yt_rsc_1_2_i_adra,
      adra_d => yt_rsc_1_2_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_2_i_da_d_1,
      qa_d => yt_rsc_1_2_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_2_i_qa <= yt_rsc_1_2_qa;
  yt_rsc_1_2_da <= yt_rsc_1_2_i_da;
  yt_rsc_1_2_adra <= yt_rsc_1_2_i_adra;
  yt_rsc_1_2_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_2_i_da_d_1 <= yt_rsc_1_2_i_da_d;
  yt_rsc_1_2_i_qa_d <= yt_rsc_1_2_i_qa_d_1;

  yt_rsc_1_3_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_42_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_3_clken,
      qa => yt_rsc_1_3_i_qa,
      wea => yt_rsc_1_3_wea,
      da => yt_rsc_1_3_i_da,
      adra => yt_rsc_1_3_i_adra,
      adra_d => yt_rsc_1_3_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_3_i_da_d_1,
      qa_d => yt_rsc_1_3_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_3_i_qa <= yt_rsc_1_3_qa;
  yt_rsc_1_3_da <= yt_rsc_1_3_i_da;
  yt_rsc_1_3_adra <= yt_rsc_1_3_i_adra;
  yt_rsc_1_3_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_3_i_da_d_1 <= yt_rsc_1_3_i_da_d;
  yt_rsc_1_3_i_qa_d <= yt_rsc_1_3_i_qa_d_1;

  yt_rsc_1_4_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_43_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_4_clken,
      qa => yt_rsc_1_4_i_qa,
      wea => yt_rsc_1_4_wea,
      da => yt_rsc_1_4_i_da,
      adra => yt_rsc_1_4_i_adra,
      adra_d => yt_rsc_1_4_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_4_i_da_d_1,
      qa_d => yt_rsc_1_4_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_4_i_qa <= yt_rsc_1_4_qa;
  yt_rsc_1_4_da <= yt_rsc_1_4_i_da;
  yt_rsc_1_4_adra <= yt_rsc_1_4_i_adra;
  yt_rsc_1_4_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_4_i_da_d_1 <= yt_rsc_1_4_i_da_d;
  yt_rsc_1_4_i_qa_d <= yt_rsc_1_4_i_qa_d_1;

  yt_rsc_1_5_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_44_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_5_clken,
      qa => yt_rsc_1_5_i_qa,
      wea => yt_rsc_1_5_wea,
      da => yt_rsc_1_5_i_da,
      adra => yt_rsc_1_5_i_adra,
      adra_d => yt_rsc_1_5_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_5_i_da_d_1,
      qa_d => yt_rsc_1_5_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_5_i_qa <= yt_rsc_1_5_qa;
  yt_rsc_1_5_da <= yt_rsc_1_5_i_da;
  yt_rsc_1_5_adra <= yt_rsc_1_5_i_adra;
  yt_rsc_1_5_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_5_i_da_d_1 <= yt_rsc_1_5_i_da_d;
  yt_rsc_1_5_i_qa_d <= yt_rsc_1_5_i_qa_d_1;

  yt_rsc_1_6_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_45_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_6_clken,
      qa => yt_rsc_1_6_i_qa,
      wea => yt_rsc_1_6_wea,
      da => yt_rsc_1_6_i_da,
      adra => yt_rsc_1_6_i_adra,
      adra_d => yt_rsc_1_6_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_6_i_da_d_1,
      qa_d => yt_rsc_1_6_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_6_i_qa <= yt_rsc_1_6_qa;
  yt_rsc_1_6_da <= yt_rsc_1_6_i_da;
  yt_rsc_1_6_adra <= yt_rsc_1_6_i_adra;
  yt_rsc_1_6_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_6_i_da_d_1 <= yt_rsc_1_6_i_da_d;
  yt_rsc_1_6_i_qa_d <= yt_rsc_1_6_i_qa_d_1;

  yt_rsc_1_7_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_46_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_7_clken,
      qa => yt_rsc_1_7_i_qa,
      wea => yt_rsc_1_7_wea,
      da => yt_rsc_1_7_i_da,
      adra => yt_rsc_1_7_i_adra,
      adra_d => yt_rsc_1_7_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_7_i_da_d_1,
      qa_d => yt_rsc_1_7_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_7_i_qa <= yt_rsc_1_7_qa;
  yt_rsc_1_7_da <= yt_rsc_1_7_i_da;
  yt_rsc_1_7_adra <= yt_rsc_1_7_i_adra;
  yt_rsc_1_7_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_7_i_da_d_1 <= yt_rsc_1_7_i_da_d;
  yt_rsc_1_7_i_qa_d <= yt_rsc_1_7_i_qa_d_1;

  yt_rsc_1_8_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_47_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_8_clken,
      qa => yt_rsc_1_8_i_qa,
      wea => yt_rsc_1_8_wea,
      da => yt_rsc_1_8_i_da,
      adra => yt_rsc_1_8_i_adra,
      adra_d => yt_rsc_1_8_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_8_i_da_d_1,
      qa_d => yt_rsc_1_8_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_8_i_qa <= yt_rsc_1_8_qa;
  yt_rsc_1_8_da <= yt_rsc_1_8_i_da;
  yt_rsc_1_8_adra <= yt_rsc_1_8_i_adra;
  yt_rsc_1_8_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_8_i_da_d_1 <= yt_rsc_1_8_i_da_d;
  yt_rsc_1_8_i_qa_d <= yt_rsc_1_8_i_qa_d_1;

  yt_rsc_1_9_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_48_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_9_clken,
      qa => yt_rsc_1_9_i_qa,
      wea => yt_rsc_1_9_wea,
      da => yt_rsc_1_9_i_da,
      adra => yt_rsc_1_9_i_adra,
      adra_d => yt_rsc_1_9_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_9_i_da_d_1,
      qa_d => yt_rsc_1_9_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_9_i_qa <= yt_rsc_1_9_qa;
  yt_rsc_1_9_da <= yt_rsc_1_9_i_da;
  yt_rsc_1_9_adra <= yt_rsc_1_9_i_adra;
  yt_rsc_1_9_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_9_i_da_d_1 <= yt_rsc_1_9_i_da_d;
  yt_rsc_1_9_i_qa_d <= yt_rsc_1_9_i_qa_d_1;

  yt_rsc_1_10_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_49_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_10_clken,
      qa => yt_rsc_1_10_i_qa,
      wea => yt_rsc_1_10_wea,
      da => yt_rsc_1_10_i_da,
      adra => yt_rsc_1_10_i_adra,
      adra_d => yt_rsc_1_10_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_10_i_da_d_1,
      qa_d => yt_rsc_1_10_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_10_i_qa <= yt_rsc_1_10_qa;
  yt_rsc_1_10_da <= yt_rsc_1_10_i_da;
  yt_rsc_1_10_adra <= yt_rsc_1_10_i_adra;
  yt_rsc_1_10_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_10_i_da_d_1 <= yt_rsc_1_10_i_da_d;
  yt_rsc_1_10_i_qa_d <= yt_rsc_1_10_i_qa_d_1;

  yt_rsc_1_11_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_50_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_11_clken,
      qa => yt_rsc_1_11_i_qa,
      wea => yt_rsc_1_11_wea,
      da => yt_rsc_1_11_i_da,
      adra => yt_rsc_1_11_i_adra,
      adra_d => yt_rsc_1_11_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_11_i_da_d_1,
      qa_d => yt_rsc_1_11_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_11_i_qa <= yt_rsc_1_11_qa;
  yt_rsc_1_11_da <= yt_rsc_1_11_i_da;
  yt_rsc_1_11_adra <= yt_rsc_1_11_i_adra;
  yt_rsc_1_11_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_11_i_da_d_1 <= yt_rsc_1_11_i_da_d;
  yt_rsc_1_11_i_qa_d <= yt_rsc_1_11_i_qa_d_1;

  yt_rsc_1_12_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_51_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_12_clken,
      qa => yt_rsc_1_12_i_qa,
      wea => yt_rsc_1_12_wea,
      da => yt_rsc_1_12_i_da,
      adra => yt_rsc_1_12_i_adra,
      adra_d => yt_rsc_1_12_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_12_i_da_d_1,
      qa_d => yt_rsc_1_12_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_12_i_qa <= yt_rsc_1_12_qa;
  yt_rsc_1_12_da <= yt_rsc_1_12_i_da;
  yt_rsc_1_12_adra <= yt_rsc_1_12_i_adra;
  yt_rsc_1_12_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_12_i_da_d_1 <= yt_rsc_1_12_i_da_d;
  yt_rsc_1_12_i_qa_d <= yt_rsc_1_12_i_qa_d_1;

  yt_rsc_1_13_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_52_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_13_clken,
      qa => yt_rsc_1_13_i_qa,
      wea => yt_rsc_1_13_wea,
      da => yt_rsc_1_13_i_da,
      adra => yt_rsc_1_13_i_adra,
      adra_d => yt_rsc_1_13_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_13_i_da_d_1,
      qa_d => yt_rsc_1_13_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_13_i_qa <= yt_rsc_1_13_qa;
  yt_rsc_1_13_da <= yt_rsc_1_13_i_da;
  yt_rsc_1_13_adra <= yt_rsc_1_13_i_adra;
  yt_rsc_1_13_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_13_i_da_d_1 <= yt_rsc_1_13_i_da_d;
  yt_rsc_1_13_i_qa_d <= yt_rsc_1_13_i_qa_d_1;

  yt_rsc_1_14_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_53_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_14_clken,
      qa => yt_rsc_1_14_i_qa,
      wea => yt_rsc_1_14_wea,
      da => yt_rsc_1_14_i_da,
      adra => yt_rsc_1_14_i_adra,
      adra_d => yt_rsc_1_14_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_14_i_da_d_1,
      qa_d => yt_rsc_1_14_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_14_i_qa <= yt_rsc_1_14_qa;
  yt_rsc_1_14_da <= yt_rsc_1_14_i_da;
  yt_rsc_1_14_adra <= yt_rsc_1_14_i_adra;
  yt_rsc_1_14_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_14_i_da_d_1 <= yt_rsc_1_14_i_da_d;
  yt_rsc_1_14_i_qa_d <= yt_rsc_1_14_i_qa_d_1;

  yt_rsc_1_15_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_54_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_15_clken,
      qa => yt_rsc_1_15_i_qa,
      wea => yt_rsc_1_15_wea,
      da => yt_rsc_1_15_i_da,
      adra => yt_rsc_1_15_i_adra,
      adra_d => yt_rsc_1_15_i_adra_d,
      clken_d => yt_rsc_1_0_i_clken_d,
      da_d => yt_rsc_1_15_i_da_d_1,
      qa_d => yt_rsc_1_15_i_qa_d_1,
      wea_d => yt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_0_i_wea_d_iff
    );
  yt_rsc_1_15_i_qa <= yt_rsc_1_15_qa;
  yt_rsc_1_15_da <= yt_rsc_1_15_i_da;
  yt_rsc_1_15_adra <= yt_rsc_1_15_i_adra;
  yt_rsc_1_15_i_adra_d <= yt_rsc_1_0_i_adra_d_iff;
  yt_rsc_1_15_i_da_d_1 <= yt_rsc_1_15_i_da_d;
  yt_rsc_1_15_i_qa_d <= yt_rsc_1_15_i_qa_d_1;

  yt_rsc_1_16_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_55_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_16_clken,
      qa => yt_rsc_1_16_i_qa,
      wea => yt_rsc_1_16_wea,
      da => yt_rsc_1_16_i_da,
      adra => yt_rsc_1_16_i_adra,
      adra_d => yt_rsc_1_16_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_16_i_da_d_1,
      qa_d => yt_rsc_1_16_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_16_i_qa <= yt_rsc_1_16_qa;
  yt_rsc_1_16_da <= yt_rsc_1_16_i_da;
  yt_rsc_1_16_adra <= yt_rsc_1_16_i_adra;
  yt_rsc_1_16_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_16_i_da_d_1 <= yt_rsc_1_16_i_da_d;
  yt_rsc_1_16_i_qa_d <= yt_rsc_1_16_i_qa_d_1;

  yt_rsc_1_17_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_56_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_17_clken,
      qa => yt_rsc_1_17_i_qa,
      wea => yt_rsc_1_17_wea,
      da => yt_rsc_1_17_i_da,
      adra => yt_rsc_1_17_i_adra,
      adra_d => yt_rsc_1_17_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_17_i_da_d_1,
      qa_d => yt_rsc_1_17_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_17_i_qa <= yt_rsc_1_17_qa;
  yt_rsc_1_17_da <= yt_rsc_1_17_i_da;
  yt_rsc_1_17_adra <= yt_rsc_1_17_i_adra;
  yt_rsc_1_17_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_17_i_da_d_1 <= yt_rsc_1_17_i_da_d;
  yt_rsc_1_17_i_qa_d <= yt_rsc_1_17_i_qa_d_1;

  yt_rsc_1_18_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_57_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_18_clken,
      qa => yt_rsc_1_18_i_qa,
      wea => yt_rsc_1_18_wea,
      da => yt_rsc_1_18_i_da,
      adra => yt_rsc_1_18_i_adra,
      adra_d => yt_rsc_1_18_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_18_i_da_d_1,
      qa_d => yt_rsc_1_18_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_18_i_qa <= yt_rsc_1_18_qa;
  yt_rsc_1_18_da <= yt_rsc_1_18_i_da;
  yt_rsc_1_18_adra <= yt_rsc_1_18_i_adra;
  yt_rsc_1_18_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_18_i_da_d_1 <= yt_rsc_1_18_i_da_d;
  yt_rsc_1_18_i_qa_d <= yt_rsc_1_18_i_qa_d_1;

  yt_rsc_1_19_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_58_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_19_clken,
      qa => yt_rsc_1_19_i_qa,
      wea => yt_rsc_1_19_wea,
      da => yt_rsc_1_19_i_da,
      adra => yt_rsc_1_19_i_adra,
      adra_d => yt_rsc_1_19_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_19_i_da_d_1,
      qa_d => yt_rsc_1_19_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_19_i_qa <= yt_rsc_1_19_qa;
  yt_rsc_1_19_da <= yt_rsc_1_19_i_da;
  yt_rsc_1_19_adra <= yt_rsc_1_19_i_adra;
  yt_rsc_1_19_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_19_i_da_d_1 <= yt_rsc_1_19_i_da_d;
  yt_rsc_1_19_i_qa_d <= yt_rsc_1_19_i_qa_d_1;

  yt_rsc_1_20_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_59_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_20_clken,
      qa => yt_rsc_1_20_i_qa,
      wea => yt_rsc_1_20_wea,
      da => yt_rsc_1_20_i_da,
      adra => yt_rsc_1_20_i_adra,
      adra_d => yt_rsc_1_20_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_20_i_da_d_1,
      qa_d => yt_rsc_1_20_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_20_i_qa <= yt_rsc_1_20_qa;
  yt_rsc_1_20_da <= yt_rsc_1_20_i_da;
  yt_rsc_1_20_adra <= yt_rsc_1_20_i_adra;
  yt_rsc_1_20_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_20_i_da_d_1 <= yt_rsc_1_20_i_da_d;
  yt_rsc_1_20_i_qa_d <= yt_rsc_1_20_i_qa_d_1;

  yt_rsc_1_21_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_60_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_21_clken,
      qa => yt_rsc_1_21_i_qa,
      wea => yt_rsc_1_21_wea,
      da => yt_rsc_1_21_i_da,
      adra => yt_rsc_1_21_i_adra,
      adra_d => yt_rsc_1_21_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_21_i_da_d_1,
      qa_d => yt_rsc_1_21_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_21_i_qa <= yt_rsc_1_21_qa;
  yt_rsc_1_21_da <= yt_rsc_1_21_i_da;
  yt_rsc_1_21_adra <= yt_rsc_1_21_i_adra;
  yt_rsc_1_21_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_21_i_da_d_1 <= yt_rsc_1_21_i_da_d;
  yt_rsc_1_21_i_qa_d <= yt_rsc_1_21_i_qa_d_1;

  yt_rsc_1_22_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_61_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_22_clken,
      qa => yt_rsc_1_22_i_qa,
      wea => yt_rsc_1_22_wea,
      da => yt_rsc_1_22_i_da,
      adra => yt_rsc_1_22_i_adra,
      adra_d => yt_rsc_1_22_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_22_i_da_d_1,
      qa_d => yt_rsc_1_22_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_22_i_qa <= yt_rsc_1_22_qa;
  yt_rsc_1_22_da <= yt_rsc_1_22_i_da;
  yt_rsc_1_22_adra <= yt_rsc_1_22_i_adra;
  yt_rsc_1_22_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_22_i_da_d_1 <= yt_rsc_1_22_i_da_d;
  yt_rsc_1_22_i_qa_d <= yt_rsc_1_22_i_qa_d_1;

  yt_rsc_1_23_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_62_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_23_clken,
      qa => yt_rsc_1_23_i_qa,
      wea => yt_rsc_1_23_wea,
      da => yt_rsc_1_23_i_da,
      adra => yt_rsc_1_23_i_adra,
      adra_d => yt_rsc_1_23_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_23_i_da_d_1,
      qa_d => yt_rsc_1_23_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_23_i_qa <= yt_rsc_1_23_qa;
  yt_rsc_1_23_da <= yt_rsc_1_23_i_da;
  yt_rsc_1_23_adra <= yt_rsc_1_23_i_adra;
  yt_rsc_1_23_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_23_i_da_d_1 <= yt_rsc_1_23_i_da_d;
  yt_rsc_1_23_i_qa_d <= yt_rsc_1_23_i_qa_d_1;

  yt_rsc_1_24_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_63_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_24_clken,
      qa => yt_rsc_1_24_i_qa,
      wea => yt_rsc_1_24_wea,
      da => yt_rsc_1_24_i_da,
      adra => yt_rsc_1_24_i_adra,
      adra_d => yt_rsc_1_24_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_24_i_da_d_1,
      qa_d => yt_rsc_1_24_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_24_i_qa <= yt_rsc_1_24_qa;
  yt_rsc_1_24_da <= yt_rsc_1_24_i_da;
  yt_rsc_1_24_adra <= yt_rsc_1_24_i_adra;
  yt_rsc_1_24_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_24_i_da_d_1 <= yt_rsc_1_24_i_da_d;
  yt_rsc_1_24_i_qa_d <= yt_rsc_1_24_i_qa_d_1;

  yt_rsc_1_25_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_64_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_25_clken,
      qa => yt_rsc_1_25_i_qa,
      wea => yt_rsc_1_25_wea,
      da => yt_rsc_1_25_i_da,
      adra => yt_rsc_1_25_i_adra,
      adra_d => yt_rsc_1_25_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_25_i_da_d_1,
      qa_d => yt_rsc_1_25_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_25_i_qa <= yt_rsc_1_25_qa;
  yt_rsc_1_25_da <= yt_rsc_1_25_i_da;
  yt_rsc_1_25_adra <= yt_rsc_1_25_i_adra;
  yt_rsc_1_25_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_25_i_da_d_1 <= yt_rsc_1_25_i_da_d;
  yt_rsc_1_25_i_qa_d <= yt_rsc_1_25_i_qa_d_1;

  yt_rsc_1_26_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_65_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_26_clken,
      qa => yt_rsc_1_26_i_qa,
      wea => yt_rsc_1_26_wea,
      da => yt_rsc_1_26_i_da,
      adra => yt_rsc_1_26_i_adra,
      adra_d => yt_rsc_1_26_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_26_i_da_d_1,
      qa_d => yt_rsc_1_26_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_26_i_qa <= yt_rsc_1_26_qa;
  yt_rsc_1_26_da <= yt_rsc_1_26_i_da;
  yt_rsc_1_26_adra <= yt_rsc_1_26_i_adra;
  yt_rsc_1_26_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_26_i_da_d_1 <= yt_rsc_1_26_i_da_d;
  yt_rsc_1_26_i_qa_d <= yt_rsc_1_26_i_qa_d_1;

  yt_rsc_1_27_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_66_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_27_clken,
      qa => yt_rsc_1_27_i_qa,
      wea => yt_rsc_1_27_wea,
      da => yt_rsc_1_27_i_da,
      adra => yt_rsc_1_27_i_adra,
      adra_d => yt_rsc_1_27_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_27_i_da_d_1,
      qa_d => yt_rsc_1_27_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_27_i_qa <= yt_rsc_1_27_qa;
  yt_rsc_1_27_da <= yt_rsc_1_27_i_da;
  yt_rsc_1_27_adra <= yt_rsc_1_27_i_adra;
  yt_rsc_1_27_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_27_i_da_d_1 <= yt_rsc_1_27_i_da_d;
  yt_rsc_1_27_i_qa_d <= yt_rsc_1_27_i_qa_d_1;

  yt_rsc_1_28_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_67_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_28_clken,
      qa => yt_rsc_1_28_i_qa,
      wea => yt_rsc_1_28_wea,
      da => yt_rsc_1_28_i_da,
      adra => yt_rsc_1_28_i_adra,
      adra_d => yt_rsc_1_28_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_28_i_da_d_1,
      qa_d => yt_rsc_1_28_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_28_i_qa <= yt_rsc_1_28_qa;
  yt_rsc_1_28_da <= yt_rsc_1_28_i_da;
  yt_rsc_1_28_adra <= yt_rsc_1_28_i_adra;
  yt_rsc_1_28_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_28_i_da_d_1 <= yt_rsc_1_28_i_da_d;
  yt_rsc_1_28_i_qa_d <= yt_rsc_1_28_i_qa_d_1;

  yt_rsc_1_29_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_68_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_29_clken,
      qa => yt_rsc_1_29_i_qa,
      wea => yt_rsc_1_29_wea,
      da => yt_rsc_1_29_i_da,
      adra => yt_rsc_1_29_i_adra,
      adra_d => yt_rsc_1_29_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_29_i_da_d_1,
      qa_d => yt_rsc_1_29_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_29_i_qa <= yt_rsc_1_29_qa;
  yt_rsc_1_29_da <= yt_rsc_1_29_i_da;
  yt_rsc_1_29_adra <= yt_rsc_1_29_i_adra;
  yt_rsc_1_29_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_29_i_da_d_1 <= yt_rsc_1_29_i_da_d;
  yt_rsc_1_29_i_qa_d <= yt_rsc_1_29_i_qa_d_1;

  yt_rsc_1_30_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_69_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_30_clken,
      qa => yt_rsc_1_30_i_qa,
      wea => yt_rsc_1_30_wea,
      da => yt_rsc_1_30_i_da,
      adra => yt_rsc_1_30_i_adra,
      adra_d => yt_rsc_1_30_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_30_i_da_d_1,
      qa_d => yt_rsc_1_30_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_30_i_qa <= yt_rsc_1_30_qa;
  yt_rsc_1_30_da <= yt_rsc_1_30_i_da;
  yt_rsc_1_30_adra <= yt_rsc_1_30_i_adra;
  yt_rsc_1_30_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_30_i_da_d_1 <= yt_rsc_1_30_i_da_d;
  yt_rsc_1_30_i_qa_d <= yt_rsc_1_30_i_qa_d_1;

  yt_rsc_1_31_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_en_70_4_32_16_16_32_1_gen
    PORT MAP(
      clken => yt_rsc_1_31_clken,
      qa => yt_rsc_1_31_i_qa,
      wea => yt_rsc_1_31_wea,
      da => yt_rsc_1_31_i_da,
      adra => yt_rsc_1_31_i_adra,
      adra_d => yt_rsc_1_31_i_adra_d,
      clken_d => yt_rsc_1_16_i_clken_d,
      da_d => yt_rsc_1_31_i_da_d_1,
      qa_d => yt_rsc_1_31_i_qa_d_1,
      wea_d => yt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      rwA_rw_ram_ir_internal_WMASK_B_d => yt_rsc_1_16_i_wea_d_iff
    );
  yt_rsc_1_31_i_qa <= yt_rsc_1_31_qa;
  yt_rsc_1_31_da <= yt_rsc_1_31_i_da;
  yt_rsc_1_31_adra <= yt_rsc_1_31_i_adra;
  yt_rsc_1_31_i_adra_d <= yt_rsc_1_16_i_adra_d_iff;
  yt_rsc_1_31_i_da_d_1 <= yt_rsc_1_31_i_da_d;
  yt_rsc_1_31_i_qa_d <= yt_rsc_1_31_i_qa_d_1;

  xt_rsc_0_0_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_71_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_0_i_qa,
      wea => xt_rsc_0_0_wea,
      da => xt_rsc_0_0_i_da,
      adra => xt_rsc_0_0_i_adra,
      adra_d => xt_rsc_0_0_i_adra_d,
      da_d => xt_rsc_0_0_i_da_d,
      qa_d => xt_rsc_0_0_i_qa_d_1,
      wea_d => xt_rsc_0_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_0_i_wea_d_iff
    );
  xt_rsc_0_0_i_qa <= xt_rsc_0_0_qa;
  xt_rsc_0_0_da <= xt_rsc_0_0_i_da;
  xt_rsc_0_0_adra <= xt_rsc_0_0_i_adra;
  xt_rsc_0_0_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_0_i_da_d <= xt_rsc_0_0_i_da_d_iff;
  xt_rsc_0_0_i_qa_d <= xt_rsc_0_0_i_qa_d_1;

  xt_rsc_0_1_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_72_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_1_i_qa,
      wea => xt_rsc_0_1_wea,
      da => xt_rsc_0_1_i_da,
      adra => xt_rsc_0_1_i_adra,
      adra_d => xt_rsc_0_1_i_adra_d,
      da_d => xt_rsc_0_1_i_da_d,
      qa_d => xt_rsc_0_1_i_qa_d_1,
      wea_d => xt_rsc_0_1_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_1_i_wea_d_iff
    );
  xt_rsc_0_1_i_qa <= xt_rsc_0_1_qa;
  xt_rsc_0_1_da <= xt_rsc_0_1_i_da;
  xt_rsc_0_1_adra <= xt_rsc_0_1_i_adra;
  xt_rsc_0_1_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_1_i_da_d <= xt_rsc_0_1_i_da_d_iff;
  xt_rsc_0_1_i_qa_d <= xt_rsc_0_1_i_qa_d_1;

  xt_rsc_0_2_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_73_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_2_i_qa,
      wea => xt_rsc_0_2_wea,
      da => xt_rsc_0_2_i_da,
      adra => xt_rsc_0_2_i_adra,
      adra_d => xt_rsc_0_2_i_adra_d,
      da_d => xt_rsc_0_2_i_da_d,
      qa_d => xt_rsc_0_2_i_qa_d_1,
      wea_d => xt_rsc_0_2_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_2_i_wea_d_iff
    );
  xt_rsc_0_2_i_qa <= xt_rsc_0_2_qa;
  xt_rsc_0_2_da <= xt_rsc_0_2_i_da;
  xt_rsc_0_2_adra <= xt_rsc_0_2_i_adra;
  xt_rsc_0_2_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_2_i_da_d <= xt_rsc_0_2_i_da_d_iff;
  xt_rsc_0_2_i_qa_d <= xt_rsc_0_2_i_qa_d_1;

  xt_rsc_0_3_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_74_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_3_i_qa,
      wea => xt_rsc_0_3_wea,
      da => xt_rsc_0_3_i_da,
      adra => xt_rsc_0_3_i_adra,
      adra_d => xt_rsc_0_3_i_adra_d,
      da_d => xt_rsc_0_3_i_da_d,
      qa_d => xt_rsc_0_3_i_qa_d_1,
      wea_d => xt_rsc_0_3_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_3_i_wea_d_iff
    );
  xt_rsc_0_3_i_qa <= xt_rsc_0_3_qa;
  xt_rsc_0_3_da <= xt_rsc_0_3_i_da;
  xt_rsc_0_3_adra <= xt_rsc_0_3_i_adra;
  xt_rsc_0_3_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_3_i_da_d <= xt_rsc_0_3_i_da_d_iff;
  xt_rsc_0_3_i_qa_d <= xt_rsc_0_3_i_qa_d_1;

  xt_rsc_0_4_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_75_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_4_i_qa,
      wea => xt_rsc_0_4_wea,
      da => xt_rsc_0_4_i_da,
      adra => xt_rsc_0_4_i_adra,
      adra_d => xt_rsc_0_4_i_adra_d,
      da_d => xt_rsc_0_4_i_da_d,
      qa_d => xt_rsc_0_4_i_qa_d_1,
      wea_d => xt_rsc_0_4_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_4_i_wea_d_iff
    );
  xt_rsc_0_4_i_qa <= xt_rsc_0_4_qa;
  xt_rsc_0_4_da <= xt_rsc_0_4_i_da;
  xt_rsc_0_4_adra <= xt_rsc_0_4_i_adra;
  xt_rsc_0_4_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_4_i_da_d <= xt_rsc_0_4_i_da_d_iff;
  xt_rsc_0_4_i_qa_d <= xt_rsc_0_4_i_qa_d_1;

  xt_rsc_0_5_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_76_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_5_i_qa,
      wea => xt_rsc_0_5_wea,
      da => xt_rsc_0_5_i_da,
      adra => xt_rsc_0_5_i_adra,
      adra_d => xt_rsc_0_5_i_adra_d,
      da_d => xt_rsc_0_5_i_da_d,
      qa_d => xt_rsc_0_5_i_qa_d_1,
      wea_d => xt_rsc_0_5_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_5_i_wea_d_iff
    );
  xt_rsc_0_5_i_qa <= xt_rsc_0_5_qa;
  xt_rsc_0_5_da <= xt_rsc_0_5_i_da;
  xt_rsc_0_5_adra <= xt_rsc_0_5_i_adra;
  xt_rsc_0_5_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_5_i_da_d <= xt_rsc_0_5_i_da_d_iff;
  xt_rsc_0_5_i_qa_d <= xt_rsc_0_5_i_qa_d_1;

  xt_rsc_0_6_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_77_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_6_i_qa,
      wea => xt_rsc_0_6_wea,
      da => xt_rsc_0_6_i_da,
      adra => xt_rsc_0_6_i_adra,
      adra_d => xt_rsc_0_6_i_adra_d,
      da_d => xt_rsc_0_6_i_da_d,
      qa_d => xt_rsc_0_6_i_qa_d_1,
      wea_d => xt_rsc_0_6_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_6_i_wea_d_iff
    );
  xt_rsc_0_6_i_qa <= xt_rsc_0_6_qa;
  xt_rsc_0_6_da <= xt_rsc_0_6_i_da;
  xt_rsc_0_6_adra <= xt_rsc_0_6_i_adra;
  xt_rsc_0_6_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_6_i_da_d <= xt_rsc_0_6_i_da_d_iff;
  xt_rsc_0_6_i_qa_d <= xt_rsc_0_6_i_qa_d_1;

  xt_rsc_0_7_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_78_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_7_i_qa,
      wea => xt_rsc_0_7_wea,
      da => xt_rsc_0_7_i_da,
      adra => xt_rsc_0_7_i_adra,
      adra_d => xt_rsc_0_7_i_adra_d,
      da_d => xt_rsc_0_7_i_da_d,
      qa_d => xt_rsc_0_7_i_qa_d_1,
      wea_d => xt_rsc_0_7_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_7_i_wea_d_iff
    );
  xt_rsc_0_7_i_qa <= xt_rsc_0_7_qa;
  xt_rsc_0_7_da <= xt_rsc_0_7_i_da;
  xt_rsc_0_7_adra <= xt_rsc_0_7_i_adra;
  xt_rsc_0_7_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_7_i_da_d <= xt_rsc_0_7_i_da_d_iff;
  xt_rsc_0_7_i_qa_d <= xt_rsc_0_7_i_qa_d_1;

  xt_rsc_0_8_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_79_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_8_i_qa,
      wea => xt_rsc_0_8_wea,
      da => xt_rsc_0_8_i_da,
      adra => xt_rsc_0_8_i_adra,
      adra_d => xt_rsc_0_8_i_adra_d,
      da_d => xt_rsc_0_8_i_da_d,
      qa_d => xt_rsc_0_8_i_qa_d_1,
      wea_d => xt_rsc_0_8_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_8_i_wea_d_iff
    );
  xt_rsc_0_8_i_qa <= xt_rsc_0_8_qa;
  xt_rsc_0_8_da <= xt_rsc_0_8_i_da;
  xt_rsc_0_8_adra <= xt_rsc_0_8_i_adra;
  xt_rsc_0_8_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_8_i_da_d <= xt_rsc_0_8_i_da_d_iff;
  xt_rsc_0_8_i_qa_d <= xt_rsc_0_8_i_qa_d_1;

  xt_rsc_0_9_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_80_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_9_i_qa,
      wea => xt_rsc_0_9_wea,
      da => xt_rsc_0_9_i_da,
      adra => xt_rsc_0_9_i_adra,
      adra_d => xt_rsc_0_9_i_adra_d,
      da_d => xt_rsc_0_9_i_da_d,
      qa_d => xt_rsc_0_9_i_qa_d_1,
      wea_d => xt_rsc_0_9_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_9_i_wea_d_iff
    );
  xt_rsc_0_9_i_qa <= xt_rsc_0_9_qa;
  xt_rsc_0_9_da <= xt_rsc_0_9_i_da;
  xt_rsc_0_9_adra <= xt_rsc_0_9_i_adra;
  xt_rsc_0_9_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_9_i_da_d <= xt_rsc_0_9_i_da_d_iff;
  xt_rsc_0_9_i_qa_d <= xt_rsc_0_9_i_qa_d_1;

  xt_rsc_0_10_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_81_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_10_i_qa,
      wea => xt_rsc_0_10_wea,
      da => xt_rsc_0_10_i_da,
      adra => xt_rsc_0_10_i_adra,
      adra_d => xt_rsc_0_10_i_adra_d,
      da_d => xt_rsc_0_10_i_da_d,
      qa_d => xt_rsc_0_10_i_qa_d_1,
      wea_d => xt_rsc_0_10_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_10_i_wea_d_iff
    );
  xt_rsc_0_10_i_qa <= xt_rsc_0_10_qa;
  xt_rsc_0_10_da <= xt_rsc_0_10_i_da;
  xt_rsc_0_10_adra <= xt_rsc_0_10_i_adra;
  xt_rsc_0_10_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_10_i_da_d <= xt_rsc_0_10_i_da_d_iff;
  xt_rsc_0_10_i_qa_d <= xt_rsc_0_10_i_qa_d_1;

  xt_rsc_0_11_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_82_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_11_i_qa,
      wea => xt_rsc_0_11_wea,
      da => xt_rsc_0_11_i_da,
      adra => xt_rsc_0_11_i_adra,
      adra_d => xt_rsc_0_11_i_adra_d,
      da_d => xt_rsc_0_11_i_da_d,
      qa_d => xt_rsc_0_11_i_qa_d_1,
      wea_d => xt_rsc_0_11_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_11_i_wea_d_iff
    );
  xt_rsc_0_11_i_qa <= xt_rsc_0_11_qa;
  xt_rsc_0_11_da <= xt_rsc_0_11_i_da;
  xt_rsc_0_11_adra <= xt_rsc_0_11_i_adra;
  xt_rsc_0_11_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_11_i_da_d <= xt_rsc_0_11_i_da_d_iff;
  xt_rsc_0_11_i_qa_d <= xt_rsc_0_11_i_qa_d_1;

  xt_rsc_0_12_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_83_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_12_i_qa,
      wea => xt_rsc_0_12_wea,
      da => xt_rsc_0_12_i_da,
      adra => xt_rsc_0_12_i_adra,
      adra_d => xt_rsc_0_12_i_adra_d,
      da_d => xt_rsc_0_12_i_da_d,
      qa_d => xt_rsc_0_12_i_qa_d_1,
      wea_d => xt_rsc_0_12_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_12_i_wea_d_iff
    );
  xt_rsc_0_12_i_qa <= xt_rsc_0_12_qa;
  xt_rsc_0_12_da <= xt_rsc_0_12_i_da;
  xt_rsc_0_12_adra <= xt_rsc_0_12_i_adra;
  xt_rsc_0_12_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_12_i_da_d <= xt_rsc_0_12_i_da_d_iff;
  xt_rsc_0_12_i_qa_d <= xt_rsc_0_12_i_qa_d_1;

  xt_rsc_0_13_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_84_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_13_i_qa,
      wea => xt_rsc_0_13_wea,
      da => xt_rsc_0_13_i_da,
      adra => xt_rsc_0_13_i_adra,
      adra_d => xt_rsc_0_13_i_adra_d,
      da_d => xt_rsc_0_13_i_da_d,
      qa_d => xt_rsc_0_13_i_qa_d_1,
      wea_d => xt_rsc_0_13_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_13_i_wea_d_iff
    );
  xt_rsc_0_13_i_qa <= xt_rsc_0_13_qa;
  xt_rsc_0_13_da <= xt_rsc_0_13_i_da;
  xt_rsc_0_13_adra <= xt_rsc_0_13_i_adra;
  xt_rsc_0_13_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_13_i_da_d <= xt_rsc_0_13_i_da_d_iff;
  xt_rsc_0_13_i_qa_d <= xt_rsc_0_13_i_qa_d_1;

  xt_rsc_0_14_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_85_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_14_i_qa,
      wea => xt_rsc_0_14_wea,
      da => xt_rsc_0_14_i_da,
      adra => xt_rsc_0_14_i_adra,
      adra_d => xt_rsc_0_14_i_adra_d,
      da_d => xt_rsc_0_14_i_da_d,
      qa_d => xt_rsc_0_14_i_qa_d_1,
      wea_d => xt_rsc_0_14_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_14_i_wea_d_iff
    );
  xt_rsc_0_14_i_qa <= xt_rsc_0_14_qa;
  xt_rsc_0_14_da <= xt_rsc_0_14_i_da;
  xt_rsc_0_14_adra <= xt_rsc_0_14_i_adra;
  xt_rsc_0_14_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_14_i_da_d <= xt_rsc_0_14_i_da_d_iff;
  xt_rsc_0_14_i_qa_d <= xt_rsc_0_14_i_qa_d_1;

  xt_rsc_0_15_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_86_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_15_i_qa,
      wea => xt_rsc_0_15_wea,
      da => xt_rsc_0_15_i_da,
      adra => xt_rsc_0_15_i_adra,
      adra_d => xt_rsc_0_15_i_adra_d,
      da_d => xt_rsc_0_15_i_da_d,
      qa_d => xt_rsc_0_15_i_qa_d_1,
      wea_d => xt_rsc_0_15_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_15_i_wea_d_iff
    );
  xt_rsc_0_15_i_qa <= xt_rsc_0_15_qa;
  xt_rsc_0_15_da <= xt_rsc_0_15_i_da;
  xt_rsc_0_15_adra <= xt_rsc_0_15_i_adra;
  xt_rsc_0_15_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_0_15_i_da_d <= xt_rsc_0_15_i_da_d_iff;
  xt_rsc_0_15_i_qa_d <= xt_rsc_0_15_i_qa_d_1;

  xt_rsc_0_16_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_87_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_16_i_qa,
      wea => xt_rsc_0_16_wea,
      da => xt_rsc_0_16_i_da,
      adra => xt_rsc_0_16_i_adra,
      adra_d => xt_rsc_0_16_i_adra_d,
      da_d => xt_rsc_0_16_i_da_d,
      qa_d => xt_rsc_0_16_i_qa_d_1,
      wea_d => xt_rsc_0_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_16_i_wea_d_iff
    );
  xt_rsc_0_16_i_qa <= xt_rsc_0_16_qa;
  xt_rsc_0_16_da <= xt_rsc_0_16_i_da;
  xt_rsc_0_16_adra <= xt_rsc_0_16_i_adra;
  xt_rsc_0_16_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_16_i_da_d <= xt_rsc_0_0_i_da_d_iff;
  xt_rsc_0_16_i_qa_d <= xt_rsc_0_16_i_qa_d_1;

  xt_rsc_0_17_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_88_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_17_i_qa,
      wea => xt_rsc_0_17_wea,
      da => xt_rsc_0_17_i_da,
      adra => xt_rsc_0_17_i_adra,
      adra_d => xt_rsc_0_17_i_adra_d,
      da_d => xt_rsc_0_17_i_da_d,
      qa_d => xt_rsc_0_17_i_qa_d_1,
      wea_d => xt_rsc_0_17_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_17_i_wea_d_iff
    );
  xt_rsc_0_17_i_qa <= xt_rsc_0_17_qa;
  xt_rsc_0_17_da <= xt_rsc_0_17_i_da;
  xt_rsc_0_17_adra <= xt_rsc_0_17_i_adra;
  xt_rsc_0_17_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_17_i_da_d <= xt_rsc_0_1_i_da_d_iff;
  xt_rsc_0_17_i_qa_d <= xt_rsc_0_17_i_qa_d_1;

  xt_rsc_0_18_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_89_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_18_i_qa,
      wea => xt_rsc_0_18_wea,
      da => xt_rsc_0_18_i_da,
      adra => xt_rsc_0_18_i_adra,
      adra_d => xt_rsc_0_18_i_adra_d,
      da_d => xt_rsc_0_18_i_da_d,
      qa_d => xt_rsc_0_18_i_qa_d_1,
      wea_d => xt_rsc_0_18_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_18_i_wea_d_iff
    );
  xt_rsc_0_18_i_qa <= xt_rsc_0_18_qa;
  xt_rsc_0_18_da <= xt_rsc_0_18_i_da;
  xt_rsc_0_18_adra <= xt_rsc_0_18_i_adra;
  xt_rsc_0_18_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_18_i_da_d <= xt_rsc_0_2_i_da_d_iff;
  xt_rsc_0_18_i_qa_d <= xt_rsc_0_18_i_qa_d_1;

  xt_rsc_0_19_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_90_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_19_i_qa,
      wea => xt_rsc_0_19_wea,
      da => xt_rsc_0_19_i_da,
      adra => xt_rsc_0_19_i_adra,
      adra_d => xt_rsc_0_19_i_adra_d,
      da_d => xt_rsc_0_19_i_da_d,
      qa_d => xt_rsc_0_19_i_qa_d_1,
      wea_d => xt_rsc_0_19_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_19_i_wea_d_iff
    );
  xt_rsc_0_19_i_qa <= xt_rsc_0_19_qa;
  xt_rsc_0_19_da <= xt_rsc_0_19_i_da;
  xt_rsc_0_19_adra <= xt_rsc_0_19_i_adra;
  xt_rsc_0_19_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_19_i_da_d <= xt_rsc_0_3_i_da_d_iff;
  xt_rsc_0_19_i_qa_d <= xt_rsc_0_19_i_qa_d_1;

  xt_rsc_0_20_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_91_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_20_i_qa,
      wea => xt_rsc_0_20_wea,
      da => xt_rsc_0_20_i_da,
      adra => xt_rsc_0_20_i_adra,
      adra_d => xt_rsc_0_20_i_adra_d,
      da_d => xt_rsc_0_20_i_da_d,
      qa_d => xt_rsc_0_20_i_qa_d_1,
      wea_d => xt_rsc_0_20_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_20_i_wea_d_iff
    );
  xt_rsc_0_20_i_qa <= xt_rsc_0_20_qa;
  xt_rsc_0_20_da <= xt_rsc_0_20_i_da;
  xt_rsc_0_20_adra <= xt_rsc_0_20_i_adra;
  xt_rsc_0_20_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_20_i_da_d <= xt_rsc_0_4_i_da_d_iff;
  xt_rsc_0_20_i_qa_d <= xt_rsc_0_20_i_qa_d_1;

  xt_rsc_0_21_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_92_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_21_i_qa,
      wea => xt_rsc_0_21_wea,
      da => xt_rsc_0_21_i_da,
      adra => xt_rsc_0_21_i_adra,
      adra_d => xt_rsc_0_21_i_adra_d,
      da_d => xt_rsc_0_21_i_da_d,
      qa_d => xt_rsc_0_21_i_qa_d_1,
      wea_d => xt_rsc_0_21_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_21_i_wea_d_iff
    );
  xt_rsc_0_21_i_qa <= xt_rsc_0_21_qa;
  xt_rsc_0_21_da <= xt_rsc_0_21_i_da;
  xt_rsc_0_21_adra <= xt_rsc_0_21_i_adra;
  xt_rsc_0_21_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_21_i_da_d <= xt_rsc_0_5_i_da_d_iff;
  xt_rsc_0_21_i_qa_d <= xt_rsc_0_21_i_qa_d_1;

  xt_rsc_0_22_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_93_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_22_i_qa,
      wea => xt_rsc_0_22_wea,
      da => xt_rsc_0_22_i_da,
      adra => xt_rsc_0_22_i_adra,
      adra_d => xt_rsc_0_22_i_adra_d,
      da_d => xt_rsc_0_22_i_da_d,
      qa_d => xt_rsc_0_22_i_qa_d_1,
      wea_d => xt_rsc_0_22_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_22_i_wea_d_iff
    );
  xt_rsc_0_22_i_qa <= xt_rsc_0_22_qa;
  xt_rsc_0_22_da <= xt_rsc_0_22_i_da;
  xt_rsc_0_22_adra <= xt_rsc_0_22_i_adra;
  xt_rsc_0_22_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_22_i_da_d <= xt_rsc_0_6_i_da_d_iff;
  xt_rsc_0_22_i_qa_d <= xt_rsc_0_22_i_qa_d_1;

  xt_rsc_0_23_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_94_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_23_i_qa,
      wea => xt_rsc_0_23_wea,
      da => xt_rsc_0_23_i_da,
      adra => xt_rsc_0_23_i_adra,
      adra_d => xt_rsc_0_23_i_adra_d,
      da_d => xt_rsc_0_23_i_da_d,
      qa_d => xt_rsc_0_23_i_qa_d_1,
      wea_d => xt_rsc_0_23_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_23_i_wea_d_iff
    );
  xt_rsc_0_23_i_qa <= xt_rsc_0_23_qa;
  xt_rsc_0_23_da <= xt_rsc_0_23_i_da;
  xt_rsc_0_23_adra <= xt_rsc_0_23_i_adra;
  xt_rsc_0_23_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_23_i_da_d <= xt_rsc_0_7_i_da_d_iff;
  xt_rsc_0_23_i_qa_d <= xt_rsc_0_23_i_qa_d_1;

  xt_rsc_0_24_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_95_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_24_i_qa,
      wea => xt_rsc_0_24_wea,
      da => xt_rsc_0_24_i_da,
      adra => xt_rsc_0_24_i_adra,
      adra_d => xt_rsc_0_24_i_adra_d,
      da_d => xt_rsc_0_24_i_da_d,
      qa_d => xt_rsc_0_24_i_qa_d_1,
      wea_d => xt_rsc_0_24_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_24_i_wea_d_iff
    );
  xt_rsc_0_24_i_qa <= xt_rsc_0_24_qa;
  xt_rsc_0_24_da <= xt_rsc_0_24_i_da;
  xt_rsc_0_24_adra <= xt_rsc_0_24_i_adra;
  xt_rsc_0_24_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_24_i_da_d <= xt_rsc_0_8_i_da_d_iff;
  xt_rsc_0_24_i_qa_d <= xt_rsc_0_24_i_qa_d_1;

  xt_rsc_0_25_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_96_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_25_i_qa,
      wea => xt_rsc_0_25_wea,
      da => xt_rsc_0_25_i_da,
      adra => xt_rsc_0_25_i_adra,
      adra_d => xt_rsc_0_25_i_adra_d,
      da_d => xt_rsc_0_25_i_da_d,
      qa_d => xt_rsc_0_25_i_qa_d_1,
      wea_d => xt_rsc_0_25_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_25_i_wea_d_iff
    );
  xt_rsc_0_25_i_qa <= xt_rsc_0_25_qa;
  xt_rsc_0_25_da <= xt_rsc_0_25_i_da;
  xt_rsc_0_25_adra <= xt_rsc_0_25_i_adra;
  xt_rsc_0_25_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_25_i_da_d <= xt_rsc_0_9_i_da_d_iff;
  xt_rsc_0_25_i_qa_d <= xt_rsc_0_25_i_qa_d_1;

  xt_rsc_0_26_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_97_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_26_i_qa,
      wea => xt_rsc_0_26_wea,
      da => xt_rsc_0_26_i_da,
      adra => xt_rsc_0_26_i_adra,
      adra_d => xt_rsc_0_26_i_adra_d,
      da_d => xt_rsc_0_26_i_da_d,
      qa_d => xt_rsc_0_26_i_qa_d_1,
      wea_d => xt_rsc_0_26_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_26_i_wea_d_iff
    );
  xt_rsc_0_26_i_qa <= xt_rsc_0_26_qa;
  xt_rsc_0_26_da <= xt_rsc_0_26_i_da;
  xt_rsc_0_26_adra <= xt_rsc_0_26_i_adra;
  xt_rsc_0_26_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_26_i_da_d <= xt_rsc_0_10_i_da_d_iff;
  xt_rsc_0_26_i_qa_d <= xt_rsc_0_26_i_qa_d_1;

  xt_rsc_0_27_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_98_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_27_i_qa,
      wea => xt_rsc_0_27_wea,
      da => xt_rsc_0_27_i_da,
      adra => xt_rsc_0_27_i_adra,
      adra_d => xt_rsc_0_27_i_adra_d,
      da_d => xt_rsc_0_27_i_da_d,
      qa_d => xt_rsc_0_27_i_qa_d_1,
      wea_d => xt_rsc_0_27_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_27_i_wea_d_iff
    );
  xt_rsc_0_27_i_qa <= xt_rsc_0_27_qa;
  xt_rsc_0_27_da <= xt_rsc_0_27_i_da;
  xt_rsc_0_27_adra <= xt_rsc_0_27_i_adra;
  xt_rsc_0_27_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_27_i_da_d <= xt_rsc_0_11_i_da_d_iff;
  xt_rsc_0_27_i_qa_d <= xt_rsc_0_27_i_qa_d_1;

  xt_rsc_0_28_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_99_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_28_i_qa,
      wea => xt_rsc_0_28_wea,
      da => xt_rsc_0_28_i_da,
      adra => xt_rsc_0_28_i_adra,
      adra_d => xt_rsc_0_28_i_adra_d,
      da_d => xt_rsc_0_28_i_da_d,
      qa_d => xt_rsc_0_28_i_qa_d_1,
      wea_d => xt_rsc_0_28_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_28_i_wea_d_iff
    );
  xt_rsc_0_28_i_qa <= xt_rsc_0_28_qa;
  xt_rsc_0_28_da <= xt_rsc_0_28_i_da;
  xt_rsc_0_28_adra <= xt_rsc_0_28_i_adra;
  xt_rsc_0_28_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_28_i_da_d <= xt_rsc_0_12_i_da_d_iff;
  xt_rsc_0_28_i_qa_d <= xt_rsc_0_28_i_qa_d_1;

  xt_rsc_0_29_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_100_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_29_i_qa,
      wea => xt_rsc_0_29_wea,
      da => xt_rsc_0_29_i_da,
      adra => xt_rsc_0_29_i_adra,
      adra_d => xt_rsc_0_29_i_adra_d,
      da_d => xt_rsc_0_29_i_da_d,
      qa_d => xt_rsc_0_29_i_qa_d_1,
      wea_d => xt_rsc_0_29_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_29_i_wea_d_iff
    );
  xt_rsc_0_29_i_qa <= xt_rsc_0_29_qa;
  xt_rsc_0_29_da <= xt_rsc_0_29_i_da;
  xt_rsc_0_29_adra <= xt_rsc_0_29_i_adra;
  xt_rsc_0_29_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_29_i_da_d <= xt_rsc_0_13_i_da_d_iff;
  xt_rsc_0_29_i_qa_d <= xt_rsc_0_29_i_qa_d_1;

  xt_rsc_0_30_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_101_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_30_i_qa,
      wea => xt_rsc_0_30_wea,
      da => xt_rsc_0_30_i_da,
      adra => xt_rsc_0_30_i_adra,
      adra_d => xt_rsc_0_30_i_adra_d,
      da_d => xt_rsc_0_30_i_da_d,
      qa_d => xt_rsc_0_30_i_qa_d_1,
      wea_d => xt_rsc_0_30_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_30_i_wea_d_iff
    );
  xt_rsc_0_30_i_qa <= xt_rsc_0_30_qa;
  xt_rsc_0_30_da <= xt_rsc_0_30_i_da;
  xt_rsc_0_30_adra <= xt_rsc_0_30_i_adra;
  xt_rsc_0_30_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_30_i_da_d <= xt_rsc_0_14_i_da_d_iff;
  xt_rsc_0_30_i_qa_d <= xt_rsc_0_30_i_qa_d_1;

  xt_rsc_0_31_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_102_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_0_31_i_qa,
      wea => xt_rsc_0_31_wea,
      da => xt_rsc_0_31_i_da,
      adra => xt_rsc_0_31_i_adra,
      adra_d => xt_rsc_0_31_i_adra_d,
      da_d => xt_rsc_0_31_i_da_d,
      qa_d => xt_rsc_0_31_i_qa_d_1,
      wea_d => xt_rsc_0_31_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_0_31_i_wea_d_iff
    );
  xt_rsc_0_31_i_qa <= xt_rsc_0_31_qa;
  xt_rsc_0_31_da <= xt_rsc_0_31_i_da;
  xt_rsc_0_31_adra <= xt_rsc_0_31_i_adra;
  xt_rsc_0_31_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_0_31_i_da_d <= xt_rsc_0_15_i_da_d_iff;
  xt_rsc_0_31_i_qa_d <= xt_rsc_0_31_i_qa_d_1;

  xt_rsc_1_0_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_103_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_0_i_qa,
      wea => xt_rsc_1_0_wea,
      da => xt_rsc_1_0_i_da,
      adra => xt_rsc_1_0_i_adra,
      adra_d => xt_rsc_1_0_i_adra_d,
      da_d => xt_rsc_1_0_i_da_d,
      qa_d => xt_rsc_1_0_i_qa_d_1,
      wea_d => xt_rsc_1_0_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_0_i_wea_d_iff
    );
  xt_rsc_1_0_i_qa <= xt_rsc_1_0_qa;
  xt_rsc_1_0_da <= xt_rsc_1_0_i_da;
  xt_rsc_1_0_adra <= xt_rsc_1_0_i_adra;
  xt_rsc_1_0_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_0_i_da_d <= xt_rsc_1_0_i_da_d_iff;
  xt_rsc_1_0_i_qa_d <= xt_rsc_1_0_i_qa_d_1;

  xt_rsc_1_1_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_104_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_1_i_qa,
      wea => xt_rsc_1_1_wea,
      da => xt_rsc_1_1_i_da,
      adra => xt_rsc_1_1_i_adra,
      adra_d => xt_rsc_1_1_i_adra_d,
      da_d => xt_rsc_1_1_i_da_d,
      qa_d => xt_rsc_1_1_i_qa_d_1,
      wea_d => xt_rsc_1_1_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_1_i_wea_d_iff
    );
  xt_rsc_1_1_i_qa <= xt_rsc_1_1_qa;
  xt_rsc_1_1_da <= xt_rsc_1_1_i_da;
  xt_rsc_1_1_adra <= xt_rsc_1_1_i_adra;
  xt_rsc_1_1_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_1_i_da_d <= xt_rsc_1_1_i_da_d_iff;
  xt_rsc_1_1_i_qa_d <= xt_rsc_1_1_i_qa_d_1;

  xt_rsc_1_2_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_105_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_2_i_qa,
      wea => xt_rsc_1_2_wea,
      da => xt_rsc_1_2_i_da,
      adra => xt_rsc_1_2_i_adra,
      adra_d => xt_rsc_1_2_i_adra_d,
      da_d => xt_rsc_1_2_i_da_d,
      qa_d => xt_rsc_1_2_i_qa_d_1,
      wea_d => xt_rsc_1_2_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_2_i_wea_d_iff
    );
  xt_rsc_1_2_i_qa <= xt_rsc_1_2_qa;
  xt_rsc_1_2_da <= xt_rsc_1_2_i_da;
  xt_rsc_1_2_adra <= xt_rsc_1_2_i_adra;
  xt_rsc_1_2_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_2_i_da_d <= xt_rsc_1_2_i_da_d_iff;
  xt_rsc_1_2_i_qa_d <= xt_rsc_1_2_i_qa_d_1;

  xt_rsc_1_3_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_106_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_3_i_qa,
      wea => xt_rsc_1_3_wea,
      da => xt_rsc_1_3_i_da,
      adra => xt_rsc_1_3_i_adra,
      adra_d => xt_rsc_1_3_i_adra_d,
      da_d => xt_rsc_1_3_i_da_d,
      qa_d => xt_rsc_1_3_i_qa_d_1,
      wea_d => xt_rsc_1_3_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_3_i_wea_d_iff
    );
  xt_rsc_1_3_i_qa <= xt_rsc_1_3_qa;
  xt_rsc_1_3_da <= xt_rsc_1_3_i_da;
  xt_rsc_1_3_adra <= xt_rsc_1_3_i_adra;
  xt_rsc_1_3_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_3_i_da_d <= xt_rsc_1_3_i_da_d_iff;
  xt_rsc_1_3_i_qa_d <= xt_rsc_1_3_i_qa_d_1;

  xt_rsc_1_4_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_107_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_4_i_qa,
      wea => xt_rsc_1_4_wea,
      da => xt_rsc_1_4_i_da,
      adra => xt_rsc_1_4_i_adra,
      adra_d => xt_rsc_1_4_i_adra_d,
      da_d => xt_rsc_1_4_i_da_d,
      qa_d => xt_rsc_1_4_i_qa_d_1,
      wea_d => xt_rsc_1_4_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_4_i_wea_d_iff
    );
  xt_rsc_1_4_i_qa <= xt_rsc_1_4_qa;
  xt_rsc_1_4_da <= xt_rsc_1_4_i_da;
  xt_rsc_1_4_adra <= xt_rsc_1_4_i_adra;
  xt_rsc_1_4_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_4_i_da_d <= xt_rsc_1_4_i_da_d_iff;
  xt_rsc_1_4_i_qa_d <= xt_rsc_1_4_i_qa_d_1;

  xt_rsc_1_5_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_108_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_5_i_qa,
      wea => xt_rsc_1_5_wea,
      da => xt_rsc_1_5_i_da,
      adra => xt_rsc_1_5_i_adra,
      adra_d => xt_rsc_1_5_i_adra_d,
      da_d => xt_rsc_1_5_i_da_d,
      qa_d => xt_rsc_1_5_i_qa_d_1,
      wea_d => xt_rsc_1_5_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_5_i_wea_d_iff
    );
  xt_rsc_1_5_i_qa <= xt_rsc_1_5_qa;
  xt_rsc_1_5_da <= xt_rsc_1_5_i_da;
  xt_rsc_1_5_adra <= xt_rsc_1_5_i_adra;
  xt_rsc_1_5_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_5_i_da_d <= xt_rsc_1_5_i_da_d_iff;
  xt_rsc_1_5_i_qa_d <= xt_rsc_1_5_i_qa_d_1;

  xt_rsc_1_6_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_109_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_6_i_qa,
      wea => xt_rsc_1_6_wea,
      da => xt_rsc_1_6_i_da,
      adra => xt_rsc_1_6_i_adra,
      adra_d => xt_rsc_1_6_i_adra_d,
      da_d => xt_rsc_1_6_i_da_d,
      qa_d => xt_rsc_1_6_i_qa_d_1,
      wea_d => xt_rsc_1_6_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_6_i_wea_d_iff
    );
  xt_rsc_1_6_i_qa <= xt_rsc_1_6_qa;
  xt_rsc_1_6_da <= xt_rsc_1_6_i_da;
  xt_rsc_1_6_adra <= xt_rsc_1_6_i_adra;
  xt_rsc_1_6_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_6_i_da_d <= xt_rsc_1_6_i_da_d_iff;
  xt_rsc_1_6_i_qa_d <= xt_rsc_1_6_i_qa_d_1;

  xt_rsc_1_7_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_110_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_7_i_qa,
      wea => xt_rsc_1_7_wea,
      da => xt_rsc_1_7_i_da,
      adra => xt_rsc_1_7_i_adra,
      adra_d => xt_rsc_1_7_i_adra_d,
      da_d => xt_rsc_1_7_i_da_d,
      qa_d => xt_rsc_1_7_i_qa_d_1,
      wea_d => xt_rsc_1_7_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_7_i_wea_d_iff
    );
  xt_rsc_1_7_i_qa <= xt_rsc_1_7_qa;
  xt_rsc_1_7_da <= xt_rsc_1_7_i_da;
  xt_rsc_1_7_adra <= xt_rsc_1_7_i_adra;
  xt_rsc_1_7_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_7_i_da_d <= xt_rsc_1_7_i_da_d_iff;
  xt_rsc_1_7_i_qa_d <= xt_rsc_1_7_i_qa_d_1;

  xt_rsc_1_8_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_111_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_8_i_qa,
      wea => xt_rsc_1_8_wea,
      da => xt_rsc_1_8_i_da,
      adra => xt_rsc_1_8_i_adra,
      adra_d => xt_rsc_1_8_i_adra_d,
      da_d => xt_rsc_1_8_i_da_d,
      qa_d => xt_rsc_1_8_i_qa_d_1,
      wea_d => xt_rsc_1_8_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_8_i_wea_d_iff
    );
  xt_rsc_1_8_i_qa <= xt_rsc_1_8_qa;
  xt_rsc_1_8_da <= xt_rsc_1_8_i_da;
  xt_rsc_1_8_adra <= xt_rsc_1_8_i_adra;
  xt_rsc_1_8_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_8_i_da_d <= xt_rsc_1_8_i_da_d_iff;
  xt_rsc_1_8_i_qa_d <= xt_rsc_1_8_i_qa_d_1;

  xt_rsc_1_9_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_112_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_9_i_qa,
      wea => xt_rsc_1_9_wea,
      da => xt_rsc_1_9_i_da,
      adra => xt_rsc_1_9_i_adra,
      adra_d => xt_rsc_1_9_i_adra_d,
      da_d => xt_rsc_1_9_i_da_d,
      qa_d => xt_rsc_1_9_i_qa_d_1,
      wea_d => xt_rsc_1_9_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_9_i_wea_d_iff
    );
  xt_rsc_1_9_i_qa <= xt_rsc_1_9_qa;
  xt_rsc_1_9_da <= xt_rsc_1_9_i_da;
  xt_rsc_1_9_adra <= xt_rsc_1_9_i_adra;
  xt_rsc_1_9_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_9_i_da_d <= xt_rsc_1_9_i_da_d_iff;
  xt_rsc_1_9_i_qa_d <= xt_rsc_1_9_i_qa_d_1;

  xt_rsc_1_10_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_113_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_10_i_qa,
      wea => xt_rsc_1_10_wea,
      da => xt_rsc_1_10_i_da,
      adra => xt_rsc_1_10_i_adra,
      adra_d => xt_rsc_1_10_i_adra_d,
      da_d => xt_rsc_1_10_i_da_d,
      qa_d => xt_rsc_1_10_i_qa_d_1,
      wea_d => xt_rsc_1_10_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_10_i_wea_d_iff
    );
  xt_rsc_1_10_i_qa <= xt_rsc_1_10_qa;
  xt_rsc_1_10_da <= xt_rsc_1_10_i_da;
  xt_rsc_1_10_adra <= xt_rsc_1_10_i_adra;
  xt_rsc_1_10_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_10_i_da_d <= xt_rsc_1_10_i_da_d_iff;
  xt_rsc_1_10_i_qa_d <= xt_rsc_1_10_i_qa_d_1;

  xt_rsc_1_11_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_114_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_11_i_qa,
      wea => xt_rsc_1_11_wea,
      da => xt_rsc_1_11_i_da,
      adra => xt_rsc_1_11_i_adra,
      adra_d => xt_rsc_1_11_i_adra_d,
      da_d => xt_rsc_1_11_i_da_d,
      qa_d => xt_rsc_1_11_i_qa_d_1,
      wea_d => xt_rsc_1_11_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_11_i_wea_d_iff
    );
  xt_rsc_1_11_i_qa <= xt_rsc_1_11_qa;
  xt_rsc_1_11_da <= xt_rsc_1_11_i_da;
  xt_rsc_1_11_adra <= xt_rsc_1_11_i_adra;
  xt_rsc_1_11_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_11_i_da_d <= xt_rsc_1_11_i_da_d_iff;
  xt_rsc_1_11_i_qa_d <= xt_rsc_1_11_i_qa_d_1;

  xt_rsc_1_12_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_115_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_12_i_qa,
      wea => xt_rsc_1_12_wea,
      da => xt_rsc_1_12_i_da,
      adra => xt_rsc_1_12_i_adra,
      adra_d => xt_rsc_1_12_i_adra_d,
      da_d => xt_rsc_1_12_i_da_d,
      qa_d => xt_rsc_1_12_i_qa_d_1,
      wea_d => xt_rsc_1_12_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_12_i_wea_d_iff
    );
  xt_rsc_1_12_i_qa <= xt_rsc_1_12_qa;
  xt_rsc_1_12_da <= xt_rsc_1_12_i_da;
  xt_rsc_1_12_adra <= xt_rsc_1_12_i_adra;
  xt_rsc_1_12_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_12_i_da_d <= xt_rsc_1_12_i_da_d_iff;
  xt_rsc_1_12_i_qa_d <= xt_rsc_1_12_i_qa_d_1;

  xt_rsc_1_13_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_116_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_13_i_qa,
      wea => xt_rsc_1_13_wea,
      da => xt_rsc_1_13_i_da,
      adra => xt_rsc_1_13_i_adra,
      adra_d => xt_rsc_1_13_i_adra_d,
      da_d => xt_rsc_1_13_i_da_d,
      qa_d => xt_rsc_1_13_i_qa_d_1,
      wea_d => xt_rsc_1_13_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_13_i_wea_d_iff
    );
  xt_rsc_1_13_i_qa <= xt_rsc_1_13_qa;
  xt_rsc_1_13_da <= xt_rsc_1_13_i_da;
  xt_rsc_1_13_adra <= xt_rsc_1_13_i_adra;
  xt_rsc_1_13_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_13_i_da_d <= xt_rsc_1_13_i_da_d_iff;
  xt_rsc_1_13_i_qa_d <= xt_rsc_1_13_i_qa_d_1;

  xt_rsc_1_14_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_117_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_14_i_qa,
      wea => xt_rsc_1_14_wea,
      da => xt_rsc_1_14_i_da,
      adra => xt_rsc_1_14_i_adra,
      adra_d => xt_rsc_1_14_i_adra_d,
      da_d => xt_rsc_1_14_i_da_d,
      qa_d => xt_rsc_1_14_i_qa_d_1,
      wea_d => xt_rsc_1_14_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_14_i_wea_d_iff
    );
  xt_rsc_1_14_i_qa <= xt_rsc_1_14_qa;
  xt_rsc_1_14_da <= xt_rsc_1_14_i_da;
  xt_rsc_1_14_adra <= xt_rsc_1_14_i_adra;
  xt_rsc_1_14_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_14_i_da_d <= xt_rsc_1_14_i_da_d_iff;
  xt_rsc_1_14_i_qa_d <= xt_rsc_1_14_i_qa_d_1;

  xt_rsc_1_15_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_118_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_15_i_qa,
      wea => xt_rsc_1_15_wea,
      da => xt_rsc_1_15_i_da,
      adra => xt_rsc_1_15_i_adra,
      adra_d => xt_rsc_1_15_i_adra_d,
      da_d => xt_rsc_1_15_i_da_d,
      qa_d => xt_rsc_1_15_i_qa_d_1,
      wea_d => xt_rsc_1_15_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_15_i_wea_d_iff
    );
  xt_rsc_1_15_i_qa <= xt_rsc_1_15_qa;
  xt_rsc_1_15_da <= xt_rsc_1_15_i_da;
  xt_rsc_1_15_adra <= xt_rsc_1_15_i_adra;
  xt_rsc_1_15_i_adra_d <= xt_rsc_0_0_i_adra_d_iff;
  xt_rsc_1_15_i_da_d <= xt_rsc_1_15_i_da_d_iff;
  xt_rsc_1_15_i_qa_d <= xt_rsc_1_15_i_qa_d_1;

  xt_rsc_1_16_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_119_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_16_i_qa,
      wea => xt_rsc_1_16_wea,
      da => xt_rsc_1_16_i_da,
      adra => xt_rsc_1_16_i_adra,
      adra_d => xt_rsc_1_16_i_adra_d,
      da_d => xt_rsc_1_16_i_da_d,
      qa_d => xt_rsc_1_16_i_qa_d_1,
      wea_d => xt_rsc_1_16_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_16_i_wea_d_iff
    );
  xt_rsc_1_16_i_qa <= xt_rsc_1_16_qa;
  xt_rsc_1_16_da <= xt_rsc_1_16_i_da;
  xt_rsc_1_16_adra <= xt_rsc_1_16_i_adra;
  xt_rsc_1_16_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_16_i_da_d <= xt_rsc_1_0_i_da_d_iff;
  xt_rsc_1_16_i_qa_d <= xt_rsc_1_16_i_qa_d_1;

  xt_rsc_1_17_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_120_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_17_i_qa,
      wea => xt_rsc_1_17_wea,
      da => xt_rsc_1_17_i_da,
      adra => xt_rsc_1_17_i_adra,
      adra_d => xt_rsc_1_17_i_adra_d,
      da_d => xt_rsc_1_17_i_da_d,
      qa_d => xt_rsc_1_17_i_qa_d_1,
      wea_d => xt_rsc_1_17_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_17_i_wea_d_iff
    );
  xt_rsc_1_17_i_qa <= xt_rsc_1_17_qa;
  xt_rsc_1_17_da <= xt_rsc_1_17_i_da;
  xt_rsc_1_17_adra <= xt_rsc_1_17_i_adra;
  xt_rsc_1_17_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_17_i_da_d <= xt_rsc_1_1_i_da_d_iff;
  xt_rsc_1_17_i_qa_d <= xt_rsc_1_17_i_qa_d_1;

  xt_rsc_1_18_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_121_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_18_i_qa,
      wea => xt_rsc_1_18_wea,
      da => xt_rsc_1_18_i_da,
      adra => xt_rsc_1_18_i_adra,
      adra_d => xt_rsc_1_18_i_adra_d,
      da_d => xt_rsc_1_18_i_da_d,
      qa_d => xt_rsc_1_18_i_qa_d_1,
      wea_d => xt_rsc_1_18_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_18_i_wea_d_iff
    );
  xt_rsc_1_18_i_qa <= xt_rsc_1_18_qa;
  xt_rsc_1_18_da <= xt_rsc_1_18_i_da;
  xt_rsc_1_18_adra <= xt_rsc_1_18_i_adra;
  xt_rsc_1_18_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_18_i_da_d <= xt_rsc_1_2_i_da_d_iff;
  xt_rsc_1_18_i_qa_d <= xt_rsc_1_18_i_qa_d_1;

  xt_rsc_1_19_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_122_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_19_i_qa,
      wea => xt_rsc_1_19_wea,
      da => xt_rsc_1_19_i_da,
      adra => xt_rsc_1_19_i_adra,
      adra_d => xt_rsc_1_19_i_adra_d,
      da_d => xt_rsc_1_19_i_da_d,
      qa_d => xt_rsc_1_19_i_qa_d_1,
      wea_d => xt_rsc_1_19_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_19_i_wea_d_iff
    );
  xt_rsc_1_19_i_qa <= xt_rsc_1_19_qa;
  xt_rsc_1_19_da <= xt_rsc_1_19_i_da;
  xt_rsc_1_19_adra <= xt_rsc_1_19_i_adra;
  xt_rsc_1_19_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_19_i_da_d <= xt_rsc_1_3_i_da_d_iff;
  xt_rsc_1_19_i_qa_d <= xt_rsc_1_19_i_qa_d_1;

  xt_rsc_1_20_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_123_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_20_i_qa,
      wea => xt_rsc_1_20_wea,
      da => xt_rsc_1_20_i_da,
      adra => xt_rsc_1_20_i_adra,
      adra_d => xt_rsc_1_20_i_adra_d,
      da_d => xt_rsc_1_20_i_da_d,
      qa_d => xt_rsc_1_20_i_qa_d_1,
      wea_d => xt_rsc_1_20_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_20_i_wea_d_iff
    );
  xt_rsc_1_20_i_qa <= xt_rsc_1_20_qa;
  xt_rsc_1_20_da <= xt_rsc_1_20_i_da;
  xt_rsc_1_20_adra <= xt_rsc_1_20_i_adra;
  xt_rsc_1_20_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_20_i_da_d <= xt_rsc_1_4_i_da_d_iff;
  xt_rsc_1_20_i_qa_d <= xt_rsc_1_20_i_qa_d_1;

  xt_rsc_1_21_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_124_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_21_i_qa,
      wea => xt_rsc_1_21_wea,
      da => xt_rsc_1_21_i_da,
      adra => xt_rsc_1_21_i_adra,
      adra_d => xt_rsc_1_21_i_adra_d,
      da_d => xt_rsc_1_21_i_da_d,
      qa_d => xt_rsc_1_21_i_qa_d_1,
      wea_d => xt_rsc_1_21_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_21_i_wea_d_iff
    );
  xt_rsc_1_21_i_qa <= xt_rsc_1_21_qa;
  xt_rsc_1_21_da <= xt_rsc_1_21_i_da;
  xt_rsc_1_21_adra <= xt_rsc_1_21_i_adra;
  xt_rsc_1_21_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_21_i_da_d <= xt_rsc_1_5_i_da_d_iff;
  xt_rsc_1_21_i_qa_d <= xt_rsc_1_21_i_qa_d_1;

  xt_rsc_1_22_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_125_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_22_i_qa,
      wea => xt_rsc_1_22_wea,
      da => xt_rsc_1_22_i_da,
      adra => xt_rsc_1_22_i_adra,
      adra_d => xt_rsc_1_22_i_adra_d,
      da_d => xt_rsc_1_22_i_da_d,
      qa_d => xt_rsc_1_22_i_qa_d_1,
      wea_d => xt_rsc_1_22_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_22_i_wea_d_iff
    );
  xt_rsc_1_22_i_qa <= xt_rsc_1_22_qa;
  xt_rsc_1_22_da <= xt_rsc_1_22_i_da;
  xt_rsc_1_22_adra <= xt_rsc_1_22_i_adra;
  xt_rsc_1_22_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_22_i_da_d <= xt_rsc_1_6_i_da_d_iff;
  xt_rsc_1_22_i_qa_d <= xt_rsc_1_22_i_qa_d_1;

  xt_rsc_1_23_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_126_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_23_i_qa,
      wea => xt_rsc_1_23_wea,
      da => xt_rsc_1_23_i_da,
      adra => xt_rsc_1_23_i_adra,
      adra_d => xt_rsc_1_23_i_adra_d,
      da_d => xt_rsc_1_23_i_da_d,
      qa_d => xt_rsc_1_23_i_qa_d_1,
      wea_d => xt_rsc_1_23_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_23_i_wea_d_iff
    );
  xt_rsc_1_23_i_qa <= xt_rsc_1_23_qa;
  xt_rsc_1_23_da <= xt_rsc_1_23_i_da;
  xt_rsc_1_23_adra <= xt_rsc_1_23_i_adra;
  xt_rsc_1_23_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_23_i_da_d <= xt_rsc_1_7_i_da_d_iff;
  xt_rsc_1_23_i_qa_d <= xt_rsc_1_23_i_qa_d_1;

  xt_rsc_1_24_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_127_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_24_i_qa,
      wea => xt_rsc_1_24_wea,
      da => xt_rsc_1_24_i_da,
      adra => xt_rsc_1_24_i_adra,
      adra_d => xt_rsc_1_24_i_adra_d,
      da_d => xt_rsc_1_24_i_da_d,
      qa_d => xt_rsc_1_24_i_qa_d_1,
      wea_d => xt_rsc_1_24_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_24_i_wea_d_iff
    );
  xt_rsc_1_24_i_qa <= xt_rsc_1_24_qa;
  xt_rsc_1_24_da <= xt_rsc_1_24_i_da;
  xt_rsc_1_24_adra <= xt_rsc_1_24_i_adra;
  xt_rsc_1_24_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_24_i_da_d <= xt_rsc_1_8_i_da_d_iff;
  xt_rsc_1_24_i_qa_d <= xt_rsc_1_24_i_qa_d_1;

  xt_rsc_1_25_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_128_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_25_i_qa,
      wea => xt_rsc_1_25_wea,
      da => xt_rsc_1_25_i_da,
      adra => xt_rsc_1_25_i_adra,
      adra_d => xt_rsc_1_25_i_adra_d,
      da_d => xt_rsc_1_25_i_da_d,
      qa_d => xt_rsc_1_25_i_qa_d_1,
      wea_d => xt_rsc_1_25_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_25_i_wea_d_iff
    );
  xt_rsc_1_25_i_qa <= xt_rsc_1_25_qa;
  xt_rsc_1_25_da <= xt_rsc_1_25_i_da;
  xt_rsc_1_25_adra <= xt_rsc_1_25_i_adra;
  xt_rsc_1_25_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_25_i_da_d <= xt_rsc_1_9_i_da_d_iff;
  xt_rsc_1_25_i_qa_d <= xt_rsc_1_25_i_qa_d_1;

  xt_rsc_1_26_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_129_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_26_i_qa,
      wea => xt_rsc_1_26_wea,
      da => xt_rsc_1_26_i_da,
      adra => xt_rsc_1_26_i_adra,
      adra_d => xt_rsc_1_26_i_adra_d,
      da_d => xt_rsc_1_26_i_da_d,
      qa_d => xt_rsc_1_26_i_qa_d_1,
      wea_d => xt_rsc_1_26_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_26_i_wea_d_iff
    );
  xt_rsc_1_26_i_qa <= xt_rsc_1_26_qa;
  xt_rsc_1_26_da <= xt_rsc_1_26_i_da;
  xt_rsc_1_26_adra <= xt_rsc_1_26_i_adra;
  xt_rsc_1_26_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_26_i_da_d <= xt_rsc_1_10_i_da_d_iff;
  xt_rsc_1_26_i_qa_d <= xt_rsc_1_26_i_qa_d_1;

  xt_rsc_1_27_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_130_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_27_i_qa,
      wea => xt_rsc_1_27_wea,
      da => xt_rsc_1_27_i_da,
      adra => xt_rsc_1_27_i_adra,
      adra_d => xt_rsc_1_27_i_adra_d,
      da_d => xt_rsc_1_27_i_da_d,
      qa_d => xt_rsc_1_27_i_qa_d_1,
      wea_d => xt_rsc_1_27_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_27_i_wea_d_iff
    );
  xt_rsc_1_27_i_qa <= xt_rsc_1_27_qa;
  xt_rsc_1_27_da <= xt_rsc_1_27_i_da;
  xt_rsc_1_27_adra <= xt_rsc_1_27_i_adra;
  xt_rsc_1_27_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_27_i_da_d <= xt_rsc_1_11_i_da_d_iff;
  xt_rsc_1_27_i_qa_d <= xt_rsc_1_27_i_qa_d_1;

  xt_rsc_1_28_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_131_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_28_i_qa,
      wea => xt_rsc_1_28_wea,
      da => xt_rsc_1_28_i_da,
      adra => xt_rsc_1_28_i_adra,
      adra_d => xt_rsc_1_28_i_adra_d,
      da_d => xt_rsc_1_28_i_da_d,
      qa_d => xt_rsc_1_28_i_qa_d_1,
      wea_d => xt_rsc_1_28_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_28_i_wea_d_iff
    );
  xt_rsc_1_28_i_qa <= xt_rsc_1_28_qa;
  xt_rsc_1_28_da <= xt_rsc_1_28_i_da;
  xt_rsc_1_28_adra <= xt_rsc_1_28_i_adra;
  xt_rsc_1_28_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_28_i_da_d <= xt_rsc_1_12_i_da_d_iff;
  xt_rsc_1_28_i_qa_d <= xt_rsc_1_28_i_qa_d_1;

  xt_rsc_1_29_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_132_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_29_i_qa,
      wea => xt_rsc_1_29_wea,
      da => xt_rsc_1_29_i_da,
      adra => xt_rsc_1_29_i_adra,
      adra_d => xt_rsc_1_29_i_adra_d,
      da_d => xt_rsc_1_29_i_da_d,
      qa_d => xt_rsc_1_29_i_qa_d_1,
      wea_d => xt_rsc_1_29_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_29_i_wea_d_iff
    );
  xt_rsc_1_29_i_qa <= xt_rsc_1_29_qa;
  xt_rsc_1_29_da <= xt_rsc_1_29_i_da;
  xt_rsc_1_29_adra <= xt_rsc_1_29_i_adra;
  xt_rsc_1_29_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_29_i_da_d <= xt_rsc_1_13_i_da_d_iff;
  xt_rsc_1_29_i_qa_d <= xt_rsc_1_29_i_qa_d_1;

  xt_rsc_1_30_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_133_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_30_i_qa,
      wea => xt_rsc_1_30_wea,
      da => xt_rsc_1_30_i_da,
      adra => xt_rsc_1_30_i_adra,
      adra_d => xt_rsc_1_30_i_adra_d,
      da_d => xt_rsc_1_30_i_da_d,
      qa_d => xt_rsc_1_30_i_qa_d_1,
      wea_d => xt_rsc_1_30_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_30_i_wea_d_iff
    );
  xt_rsc_1_30_i_qa <= xt_rsc_1_30_qa;
  xt_rsc_1_30_da <= xt_rsc_1_30_i_da;
  xt_rsc_1_30_adra <= xt_rsc_1_30_i_adra;
  xt_rsc_1_30_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_30_i_da_d <= xt_rsc_1_14_i_da_d_iff;
  xt_rsc_1_30_i_qa_d <= xt_rsc_1_30_i_qa_d_1;

  xt_rsc_1_31_i : peaseNTT_Xilinx_RAMS_BLOCK_2R1W_RBW_rwport_134_4_32_16_16_32_1_gen
    PORT MAP(
      qa => xt_rsc_1_31_i_qa,
      wea => xt_rsc_1_31_wea,
      da => xt_rsc_1_31_i_da,
      adra => xt_rsc_1_31_i_adra,
      adra_d => xt_rsc_1_31_i_adra_d,
      da_d => xt_rsc_1_31_i_da_d,
      qa_d => xt_rsc_1_31_i_qa_d_1,
      wea_d => xt_rsc_1_31_i_wea_d_iff,
      rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      rwA_rw_ram_ir_internal_WMASK_B_d => xt_rsc_1_31_i_wea_d_iff
    );
  xt_rsc_1_31_i_qa <= xt_rsc_1_31_qa;
  xt_rsc_1_31_da <= xt_rsc_1_31_i_da;
  xt_rsc_1_31_adra <= xt_rsc_1_31_i_adra;
  xt_rsc_1_31_i_adra_d <= xt_rsc_0_16_i_adra_d_iff;
  xt_rsc_1_31_i_da_d <= xt_rsc_1_15_i_da_d_iff;
  xt_rsc_1_31_i_qa_d <= xt_rsc_1_31_i_qa_d_1;

  peaseNTT_core_inst : peaseNTT_core
    PORT MAP(
      clk => clk,
      rst => rst,
      xt_rsc_triosy_0_0_lz => xt_rsc_triosy_0_0_lz,
      xt_rsc_triosy_0_1_lz => xt_rsc_triosy_0_1_lz,
      xt_rsc_triosy_0_2_lz => xt_rsc_triosy_0_2_lz,
      xt_rsc_triosy_0_3_lz => xt_rsc_triosy_0_3_lz,
      xt_rsc_triosy_0_4_lz => xt_rsc_triosy_0_4_lz,
      xt_rsc_triosy_0_5_lz => xt_rsc_triosy_0_5_lz,
      xt_rsc_triosy_0_6_lz => xt_rsc_triosy_0_6_lz,
      xt_rsc_triosy_0_7_lz => xt_rsc_triosy_0_7_lz,
      xt_rsc_triosy_0_8_lz => xt_rsc_triosy_0_8_lz,
      xt_rsc_triosy_0_9_lz => xt_rsc_triosy_0_9_lz,
      xt_rsc_triosy_0_10_lz => xt_rsc_triosy_0_10_lz,
      xt_rsc_triosy_0_11_lz => xt_rsc_triosy_0_11_lz,
      xt_rsc_triosy_0_12_lz => xt_rsc_triosy_0_12_lz,
      xt_rsc_triosy_0_13_lz => xt_rsc_triosy_0_13_lz,
      xt_rsc_triosy_0_14_lz => xt_rsc_triosy_0_14_lz,
      xt_rsc_triosy_0_15_lz => xt_rsc_triosy_0_15_lz,
      xt_rsc_triosy_0_16_lz => xt_rsc_triosy_0_16_lz,
      xt_rsc_triosy_0_17_lz => xt_rsc_triosy_0_17_lz,
      xt_rsc_triosy_0_18_lz => xt_rsc_triosy_0_18_lz,
      xt_rsc_triosy_0_19_lz => xt_rsc_triosy_0_19_lz,
      xt_rsc_triosy_0_20_lz => xt_rsc_triosy_0_20_lz,
      xt_rsc_triosy_0_21_lz => xt_rsc_triosy_0_21_lz,
      xt_rsc_triosy_0_22_lz => xt_rsc_triosy_0_22_lz,
      xt_rsc_triosy_0_23_lz => xt_rsc_triosy_0_23_lz,
      xt_rsc_triosy_0_24_lz => xt_rsc_triosy_0_24_lz,
      xt_rsc_triosy_0_25_lz => xt_rsc_triosy_0_25_lz,
      xt_rsc_triosy_0_26_lz => xt_rsc_triosy_0_26_lz,
      xt_rsc_triosy_0_27_lz => xt_rsc_triosy_0_27_lz,
      xt_rsc_triosy_0_28_lz => xt_rsc_triosy_0_28_lz,
      xt_rsc_triosy_0_29_lz => xt_rsc_triosy_0_29_lz,
      xt_rsc_triosy_0_30_lz => xt_rsc_triosy_0_30_lz,
      xt_rsc_triosy_0_31_lz => xt_rsc_triosy_0_31_lz,
      xt_rsc_triosy_1_0_lz => xt_rsc_triosy_1_0_lz,
      xt_rsc_triosy_1_1_lz => xt_rsc_triosy_1_1_lz,
      xt_rsc_triosy_1_2_lz => xt_rsc_triosy_1_2_lz,
      xt_rsc_triosy_1_3_lz => xt_rsc_triosy_1_3_lz,
      xt_rsc_triosy_1_4_lz => xt_rsc_triosy_1_4_lz,
      xt_rsc_triosy_1_5_lz => xt_rsc_triosy_1_5_lz,
      xt_rsc_triosy_1_6_lz => xt_rsc_triosy_1_6_lz,
      xt_rsc_triosy_1_7_lz => xt_rsc_triosy_1_7_lz,
      xt_rsc_triosy_1_8_lz => xt_rsc_triosy_1_8_lz,
      xt_rsc_triosy_1_9_lz => xt_rsc_triosy_1_9_lz,
      xt_rsc_triosy_1_10_lz => xt_rsc_triosy_1_10_lz,
      xt_rsc_triosy_1_11_lz => xt_rsc_triosy_1_11_lz,
      xt_rsc_triosy_1_12_lz => xt_rsc_triosy_1_12_lz,
      xt_rsc_triosy_1_13_lz => xt_rsc_triosy_1_13_lz,
      xt_rsc_triosy_1_14_lz => xt_rsc_triosy_1_14_lz,
      xt_rsc_triosy_1_15_lz => xt_rsc_triosy_1_15_lz,
      xt_rsc_triosy_1_16_lz => xt_rsc_triosy_1_16_lz,
      xt_rsc_triosy_1_17_lz => xt_rsc_triosy_1_17_lz,
      xt_rsc_triosy_1_18_lz => xt_rsc_triosy_1_18_lz,
      xt_rsc_triosy_1_19_lz => xt_rsc_triosy_1_19_lz,
      xt_rsc_triosy_1_20_lz => xt_rsc_triosy_1_20_lz,
      xt_rsc_triosy_1_21_lz => xt_rsc_triosy_1_21_lz,
      xt_rsc_triosy_1_22_lz => xt_rsc_triosy_1_22_lz,
      xt_rsc_triosy_1_23_lz => xt_rsc_triosy_1_23_lz,
      xt_rsc_triosy_1_24_lz => xt_rsc_triosy_1_24_lz,
      xt_rsc_triosy_1_25_lz => xt_rsc_triosy_1_25_lz,
      xt_rsc_triosy_1_26_lz => xt_rsc_triosy_1_26_lz,
      xt_rsc_triosy_1_27_lz => xt_rsc_triosy_1_27_lz,
      xt_rsc_triosy_1_28_lz => xt_rsc_triosy_1_28_lz,
      xt_rsc_triosy_1_29_lz => xt_rsc_triosy_1_29_lz,
      xt_rsc_triosy_1_30_lz => xt_rsc_triosy_1_30_lz,
      xt_rsc_triosy_1_31_lz => xt_rsc_triosy_1_31_lz,
      p_rsc_dat => peaseNTT_core_inst_p_rsc_dat,
      p_rsc_triosy_lz => p_rsc_triosy_lz,
      r_rsc_triosy_lz => r_rsc_triosy_lz,
      twiddle_rsc_0_0_s_tdone => twiddle_rsc_0_0_s_tdone,
      twiddle_rsc_0_0_tr_write_done => twiddle_rsc_0_0_tr_write_done,
      twiddle_rsc_0_0_RREADY => twiddle_rsc_0_0_RREADY,
      twiddle_rsc_0_0_RVALID => twiddle_rsc_0_0_RVALID,
      twiddle_rsc_0_0_RUSER => twiddle_rsc_0_0_RUSER,
      twiddle_rsc_0_0_RLAST => twiddle_rsc_0_0_RLAST,
      twiddle_rsc_0_0_RRESP => peaseNTT_core_inst_twiddle_rsc_0_0_RRESP,
      twiddle_rsc_0_0_RDATA => peaseNTT_core_inst_twiddle_rsc_0_0_RDATA,
      twiddle_rsc_0_0_RID => twiddle_rsc_0_0_RID,
      twiddle_rsc_0_0_ARREADY => twiddle_rsc_0_0_ARREADY,
      twiddle_rsc_0_0_ARVALID => twiddle_rsc_0_0_ARVALID,
      twiddle_rsc_0_0_ARUSER => twiddle_rsc_0_0_ARUSER,
      twiddle_rsc_0_0_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_0_ARREGION,
      twiddle_rsc_0_0_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_0_ARQOS,
      twiddle_rsc_0_0_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_0_ARPROT,
      twiddle_rsc_0_0_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_0_ARCACHE,
      twiddle_rsc_0_0_ARLOCK => twiddle_rsc_0_0_ARLOCK,
      twiddle_rsc_0_0_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_0_ARBURST,
      twiddle_rsc_0_0_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_0_ARSIZE,
      twiddle_rsc_0_0_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_0_ARLEN,
      twiddle_rsc_0_0_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_0_ARADDR,
      twiddle_rsc_0_0_ARID => twiddle_rsc_0_0_ARID,
      twiddle_rsc_0_0_BREADY => twiddle_rsc_0_0_BREADY,
      twiddle_rsc_0_0_BVALID => twiddle_rsc_0_0_BVALID,
      twiddle_rsc_0_0_BUSER => twiddle_rsc_0_0_BUSER,
      twiddle_rsc_0_0_BRESP => peaseNTT_core_inst_twiddle_rsc_0_0_BRESP,
      twiddle_rsc_0_0_BID => twiddle_rsc_0_0_BID,
      twiddle_rsc_0_0_WREADY => twiddle_rsc_0_0_WREADY,
      twiddle_rsc_0_0_WVALID => twiddle_rsc_0_0_WVALID,
      twiddle_rsc_0_0_WUSER => twiddle_rsc_0_0_WUSER,
      twiddle_rsc_0_0_WLAST => twiddle_rsc_0_0_WLAST,
      twiddle_rsc_0_0_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_0_WSTRB,
      twiddle_rsc_0_0_WDATA => peaseNTT_core_inst_twiddle_rsc_0_0_WDATA,
      twiddle_rsc_0_0_AWREADY => twiddle_rsc_0_0_AWREADY,
      twiddle_rsc_0_0_AWVALID => twiddle_rsc_0_0_AWVALID,
      twiddle_rsc_0_0_AWUSER => twiddle_rsc_0_0_AWUSER,
      twiddle_rsc_0_0_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_0_AWREGION,
      twiddle_rsc_0_0_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_0_AWQOS,
      twiddle_rsc_0_0_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_0_AWPROT,
      twiddle_rsc_0_0_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_0_AWCACHE,
      twiddle_rsc_0_0_AWLOCK => twiddle_rsc_0_0_AWLOCK,
      twiddle_rsc_0_0_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_0_AWBURST,
      twiddle_rsc_0_0_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_0_AWSIZE,
      twiddle_rsc_0_0_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_0_AWLEN,
      twiddle_rsc_0_0_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_0_AWADDR,
      twiddle_rsc_0_0_AWID => twiddle_rsc_0_0_AWID,
      twiddle_rsc_triosy_0_0_lz => twiddle_rsc_triosy_0_0_lz,
      twiddle_rsc_0_1_s_tdone => twiddle_rsc_0_1_s_tdone,
      twiddle_rsc_0_1_tr_write_done => twiddle_rsc_0_1_tr_write_done,
      twiddle_rsc_0_1_RREADY => twiddle_rsc_0_1_RREADY,
      twiddle_rsc_0_1_RVALID => twiddle_rsc_0_1_RVALID,
      twiddle_rsc_0_1_RUSER => twiddle_rsc_0_1_RUSER,
      twiddle_rsc_0_1_RLAST => twiddle_rsc_0_1_RLAST,
      twiddle_rsc_0_1_RRESP => peaseNTT_core_inst_twiddle_rsc_0_1_RRESP,
      twiddle_rsc_0_1_RDATA => peaseNTT_core_inst_twiddle_rsc_0_1_RDATA,
      twiddle_rsc_0_1_RID => twiddle_rsc_0_1_RID,
      twiddle_rsc_0_1_ARREADY => twiddle_rsc_0_1_ARREADY,
      twiddle_rsc_0_1_ARVALID => twiddle_rsc_0_1_ARVALID,
      twiddle_rsc_0_1_ARUSER => twiddle_rsc_0_1_ARUSER,
      twiddle_rsc_0_1_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_1_ARREGION,
      twiddle_rsc_0_1_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_1_ARQOS,
      twiddle_rsc_0_1_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_1_ARPROT,
      twiddle_rsc_0_1_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_1_ARCACHE,
      twiddle_rsc_0_1_ARLOCK => twiddle_rsc_0_1_ARLOCK,
      twiddle_rsc_0_1_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_1_ARBURST,
      twiddle_rsc_0_1_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_1_ARSIZE,
      twiddle_rsc_0_1_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_1_ARLEN,
      twiddle_rsc_0_1_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_1_ARADDR,
      twiddle_rsc_0_1_ARID => twiddle_rsc_0_1_ARID,
      twiddle_rsc_0_1_BREADY => twiddle_rsc_0_1_BREADY,
      twiddle_rsc_0_1_BVALID => twiddle_rsc_0_1_BVALID,
      twiddle_rsc_0_1_BUSER => twiddle_rsc_0_1_BUSER,
      twiddle_rsc_0_1_BRESP => peaseNTT_core_inst_twiddle_rsc_0_1_BRESP,
      twiddle_rsc_0_1_BID => twiddle_rsc_0_1_BID,
      twiddle_rsc_0_1_WREADY => twiddle_rsc_0_1_WREADY,
      twiddle_rsc_0_1_WVALID => twiddle_rsc_0_1_WVALID,
      twiddle_rsc_0_1_WUSER => twiddle_rsc_0_1_WUSER,
      twiddle_rsc_0_1_WLAST => twiddle_rsc_0_1_WLAST,
      twiddle_rsc_0_1_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_1_WSTRB,
      twiddle_rsc_0_1_WDATA => peaseNTT_core_inst_twiddle_rsc_0_1_WDATA,
      twiddle_rsc_0_1_AWREADY => twiddle_rsc_0_1_AWREADY,
      twiddle_rsc_0_1_AWVALID => twiddle_rsc_0_1_AWVALID,
      twiddle_rsc_0_1_AWUSER => twiddle_rsc_0_1_AWUSER,
      twiddle_rsc_0_1_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_1_AWREGION,
      twiddle_rsc_0_1_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_1_AWQOS,
      twiddle_rsc_0_1_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_1_AWPROT,
      twiddle_rsc_0_1_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_1_AWCACHE,
      twiddle_rsc_0_1_AWLOCK => twiddle_rsc_0_1_AWLOCK,
      twiddle_rsc_0_1_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_1_AWBURST,
      twiddle_rsc_0_1_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_1_AWSIZE,
      twiddle_rsc_0_1_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_1_AWLEN,
      twiddle_rsc_0_1_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_1_AWADDR,
      twiddle_rsc_0_1_AWID => twiddle_rsc_0_1_AWID,
      twiddle_rsc_triosy_0_1_lz => twiddle_rsc_triosy_0_1_lz,
      twiddle_rsc_0_2_s_tdone => twiddle_rsc_0_2_s_tdone,
      twiddle_rsc_0_2_tr_write_done => twiddle_rsc_0_2_tr_write_done,
      twiddle_rsc_0_2_RREADY => twiddle_rsc_0_2_RREADY,
      twiddle_rsc_0_2_RVALID => twiddle_rsc_0_2_RVALID,
      twiddle_rsc_0_2_RUSER => twiddle_rsc_0_2_RUSER,
      twiddle_rsc_0_2_RLAST => twiddle_rsc_0_2_RLAST,
      twiddle_rsc_0_2_RRESP => peaseNTT_core_inst_twiddle_rsc_0_2_RRESP,
      twiddle_rsc_0_2_RDATA => peaseNTT_core_inst_twiddle_rsc_0_2_RDATA,
      twiddle_rsc_0_2_RID => twiddle_rsc_0_2_RID,
      twiddle_rsc_0_2_ARREADY => twiddle_rsc_0_2_ARREADY,
      twiddle_rsc_0_2_ARVALID => twiddle_rsc_0_2_ARVALID,
      twiddle_rsc_0_2_ARUSER => twiddle_rsc_0_2_ARUSER,
      twiddle_rsc_0_2_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_2_ARREGION,
      twiddle_rsc_0_2_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_2_ARQOS,
      twiddle_rsc_0_2_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_2_ARPROT,
      twiddle_rsc_0_2_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_2_ARCACHE,
      twiddle_rsc_0_2_ARLOCK => twiddle_rsc_0_2_ARLOCK,
      twiddle_rsc_0_2_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_2_ARBURST,
      twiddle_rsc_0_2_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_2_ARSIZE,
      twiddle_rsc_0_2_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_2_ARLEN,
      twiddle_rsc_0_2_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_2_ARADDR,
      twiddle_rsc_0_2_ARID => twiddle_rsc_0_2_ARID,
      twiddle_rsc_0_2_BREADY => twiddle_rsc_0_2_BREADY,
      twiddle_rsc_0_2_BVALID => twiddle_rsc_0_2_BVALID,
      twiddle_rsc_0_2_BUSER => twiddle_rsc_0_2_BUSER,
      twiddle_rsc_0_2_BRESP => peaseNTT_core_inst_twiddle_rsc_0_2_BRESP,
      twiddle_rsc_0_2_BID => twiddle_rsc_0_2_BID,
      twiddle_rsc_0_2_WREADY => twiddle_rsc_0_2_WREADY,
      twiddle_rsc_0_2_WVALID => twiddle_rsc_0_2_WVALID,
      twiddle_rsc_0_2_WUSER => twiddle_rsc_0_2_WUSER,
      twiddle_rsc_0_2_WLAST => twiddle_rsc_0_2_WLAST,
      twiddle_rsc_0_2_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_2_WSTRB,
      twiddle_rsc_0_2_WDATA => peaseNTT_core_inst_twiddle_rsc_0_2_WDATA,
      twiddle_rsc_0_2_AWREADY => twiddle_rsc_0_2_AWREADY,
      twiddle_rsc_0_2_AWVALID => twiddle_rsc_0_2_AWVALID,
      twiddle_rsc_0_2_AWUSER => twiddle_rsc_0_2_AWUSER,
      twiddle_rsc_0_2_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_2_AWREGION,
      twiddle_rsc_0_2_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_2_AWQOS,
      twiddle_rsc_0_2_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_2_AWPROT,
      twiddle_rsc_0_2_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_2_AWCACHE,
      twiddle_rsc_0_2_AWLOCK => twiddle_rsc_0_2_AWLOCK,
      twiddle_rsc_0_2_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_2_AWBURST,
      twiddle_rsc_0_2_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_2_AWSIZE,
      twiddle_rsc_0_2_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_2_AWLEN,
      twiddle_rsc_0_2_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_2_AWADDR,
      twiddle_rsc_0_2_AWID => twiddle_rsc_0_2_AWID,
      twiddle_rsc_triosy_0_2_lz => twiddle_rsc_triosy_0_2_lz,
      twiddle_rsc_0_3_s_tdone => twiddle_rsc_0_3_s_tdone,
      twiddle_rsc_0_3_tr_write_done => twiddle_rsc_0_3_tr_write_done,
      twiddle_rsc_0_3_RREADY => twiddle_rsc_0_3_RREADY,
      twiddle_rsc_0_3_RVALID => twiddle_rsc_0_3_RVALID,
      twiddle_rsc_0_3_RUSER => twiddle_rsc_0_3_RUSER,
      twiddle_rsc_0_3_RLAST => twiddle_rsc_0_3_RLAST,
      twiddle_rsc_0_3_RRESP => peaseNTT_core_inst_twiddle_rsc_0_3_RRESP,
      twiddle_rsc_0_3_RDATA => peaseNTT_core_inst_twiddle_rsc_0_3_RDATA,
      twiddle_rsc_0_3_RID => twiddle_rsc_0_3_RID,
      twiddle_rsc_0_3_ARREADY => twiddle_rsc_0_3_ARREADY,
      twiddle_rsc_0_3_ARVALID => twiddle_rsc_0_3_ARVALID,
      twiddle_rsc_0_3_ARUSER => twiddle_rsc_0_3_ARUSER,
      twiddle_rsc_0_3_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_3_ARREGION,
      twiddle_rsc_0_3_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_3_ARQOS,
      twiddle_rsc_0_3_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_3_ARPROT,
      twiddle_rsc_0_3_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_3_ARCACHE,
      twiddle_rsc_0_3_ARLOCK => twiddle_rsc_0_3_ARLOCK,
      twiddle_rsc_0_3_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_3_ARBURST,
      twiddle_rsc_0_3_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_3_ARSIZE,
      twiddle_rsc_0_3_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_3_ARLEN,
      twiddle_rsc_0_3_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_3_ARADDR,
      twiddle_rsc_0_3_ARID => twiddle_rsc_0_3_ARID,
      twiddle_rsc_0_3_BREADY => twiddle_rsc_0_3_BREADY,
      twiddle_rsc_0_3_BVALID => twiddle_rsc_0_3_BVALID,
      twiddle_rsc_0_3_BUSER => twiddle_rsc_0_3_BUSER,
      twiddle_rsc_0_3_BRESP => peaseNTT_core_inst_twiddle_rsc_0_3_BRESP,
      twiddle_rsc_0_3_BID => twiddle_rsc_0_3_BID,
      twiddle_rsc_0_3_WREADY => twiddle_rsc_0_3_WREADY,
      twiddle_rsc_0_3_WVALID => twiddle_rsc_0_3_WVALID,
      twiddle_rsc_0_3_WUSER => twiddle_rsc_0_3_WUSER,
      twiddle_rsc_0_3_WLAST => twiddle_rsc_0_3_WLAST,
      twiddle_rsc_0_3_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_3_WSTRB,
      twiddle_rsc_0_3_WDATA => peaseNTT_core_inst_twiddle_rsc_0_3_WDATA,
      twiddle_rsc_0_3_AWREADY => twiddle_rsc_0_3_AWREADY,
      twiddle_rsc_0_3_AWVALID => twiddle_rsc_0_3_AWVALID,
      twiddle_rsc_0_3_AWUSER => twiddle_rsc_0_3_AWUSER,
      twiddle_rsc_0_3_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_3_AWREGION,
      twiddle_rsc_0_3_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_3_AWQOS,
      twiddle_rsc_0_3_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_3_AWPROT,
      twiddle_rsc_0_3_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_3_AWCACHE,
      twiddle_rsc_0_3_AWLOCK => twiddle_rsc_0_3_AWLOCK,
      twiddle_rsc_0_3_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_3_AWBURST,
      twiddle_rsc_0_3_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_3_AWSIZE,
      twiddle_rsc_0_3_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_3_AWLEN,
      twiddle_rsc_0_3_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_3_AWADDR,
      twiddle_rsc_0_3_AWID => twiddle_rsc_0_3_AWID,
      twiddle_rsc_triosy_0_3_lz => twiddle_rsc_triosy_0_3_lz,
      twiddle_rsc_0_4_s_tdone => twiddle_rsc_0_4_s_tdone,
      twiddle_rsc_0_4_tr_write_done => twiddle_rsc_0_4_tr_write_done,
      twiddle_rsc_0_4_RREADY => twiddle_rsc_0_4_RREADY,
      twiddle_rsc_0_4_RVALID => twiddle_rsc_0_4_RVALID,
      twiddle_rsc_0_4_RUSER => twiddle_rsc_0_4_RUSER,
      twiddle_rsc_0_4_RLAST => twiddle_rsc_0_4_RLAST,
      twiddle_rsc_0_4_RRESP => peaseNTT_core_inst_twiddle_rsc_0_4_RRESP,
      twiddle_rsc_0_4_RDATA => peaseNTT_core_inst_twiddle_rsc_0_4_RDATA,
      twiddle_rsc_0_4_RID => twiddle_rsc_0_4_RID,
      twiddle_rsc_0_4_ARREADY => twiddle_rsc_0_4_ARREADY,
      twiddle_rsc_0_4_ARVALID => twiddle_rsc_0_4_ARVALID,
      twiddle_rsc_0_4_ARUSER => twiddle_rsc_0_4_ARUSER,
      twiddle_rsc_0_4_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_4_ARREGION,
      twiddle_rsc_0_4_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_4_ARQOS,
      twiddle_rsc_0_4_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_4_ARPROT,
      twiddle_rsc_0_4_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_4_ARCACHE,
      twiddle_rsc_0_4_ARLOCK => twiddle_rsc_0_4_ARLOCK,
      twiddle_rsc_0_4_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_4_ARBURST,
      twiddle_rsc_0_4_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_4_ARSIZE,
      twiddle_rsc_0_4_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_4_ARLEN,
      twiddle_rsc_0_4_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_4_ARADDR,
      twiddle_rsc_0_4_ARID => twiddle_rsc_0_4_ARID,
      twiddle_rsc_0_4_BREADY => twiddle_rsc_0_4_BREADY,
      twiddle_rsc_0_4_BVALID => twiddle_rsc_0_4_BVALID,
      twiddle_rsc_0_4_BUSER => twiddle_rsc_0_4_BUSER,
      twiddle_rsc_0_4_BRESP => peaseNTT_core_inst_twiddle_rsc_0_4_BRESP,
      twiddle_rsc_0_4_BID => twiddle_rsc_0_4_BID,
      twiddle_rsc_0_4_WREADY => twiddle_rsc_0_4_WREADY,
      twiddle_rsc_0_4_WVALID => twiddle_rsc_0_4_WVALID,
      twiddle_rsc_0_4_WUSER => twiddle_rsc_0_4_WUSER,
      twiddle_rsc_0_4_WLAST => twiddle_rsc_0_4_WLAST,
      twiddle_rsc_0_4_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_4_WSTRB,
      twiddle_rsc_0_4_WDATA => peaseNTT_core_inst_twiddle_rsc_0_4_WDATA,
      twiddle_rsc_0_4_AWREADY => twiddle_rsc_0_4_AWREADY,
      twiddle_rsc_0_4_AWVALID => twiddle_rsc_0_4_AWVALID,
      twiddle_rsc_0_4_AWUSER => twiddle_rsc_0_4_AWUSER,
      twiddle_rsc_0_4_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_4_AWREGION,
      twiddle_rsc_0_4_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_4_AWQOS,
      twiddle_rsc_0_4_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_4_AWPROT,
      twiddle_rsc_0_4_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_4_AWCACHE,
      twiddle_rsc_0_4_AWLOCK => twiddle_rsc_0_4_AWLOCK,
      twiddle_rsc_0_4_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_4_AWBURST,
      twiddle_rsc_0_4_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_4_AWSIZE,
      twiddle_rsc_0_4_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_4_AWLEN,
      twiddle_rsc_0_4_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_4_AWADDR,
      twiddle_rsc_0_4_AWID => twiddle_rsc_0_4_AWID,
      twiddle_rsc_triosy_0_4_lz => twiddle_rsc_triosy_0_4_lz,
      twiddle_rsc_0_5_s_tdone => twiddle_rsc_0_5_s_tdone,
      twiddle_rsc_0_5_tr_write_done => twiddle_rsc_0_5_tr_write_done,
      twiddle_rsc_0_5_RREADY => twiddle_rsc_0_5_RREADY,
      twiddle_rsc_0_5_RVALID => twiddle_rsc_0_5_RVALID,
      twiddle_rsc_0_5_RUSER => twiddle_rsc_0_5_RUSER,
      twiddle_rsc_0_5_RLAST => twiddle_rsc_0_5_RLAST,
      twiddle_rsc_0_5_RRESP => peaseNTT_core_inst_twiddle_rsc_0_5_RRESP,
      twiddle_rsc_0_5_RDATA => peaseNTT_core_inst_twiddle_rsc_0_5_RDATA,
      twiddle_rsc_0_5_RID => twiddle_rsc_0_5_RID,
      twiddle_rsc_0_5_ARREADY => twiddle_rsc_0_5_ARREADY,
      twiddle_rsc_0_5_ARVALID => twiddle_rsc_0_5_ARVALID,
      twiddle_rsc_0_5_ARUSER => twiddle_rsc_0_5_ARUSER,
      twiddle_rsc_0_5_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_5_ARREGION,
      twiddle_rsc_0_5_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_5_ARQOS,
      twiddle_rsc_0_5_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_5_ARPROT,
      twiddle_rsc_0_5_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_5_ARCACHE,
      twiddle_rsc_0_5_ARLOCK => twiddle_rsc_0_5_ARLOCK,
      twiddle_rsc_0_5_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_5_ARBURST,
      twiddle_rsc_0_5_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_5_ARSIZE,
      twiddle_rsc_0_5_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_5_ARLEN,
      twiddle_rsc_0_5_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_5_ARADDR,
      twiddle_rsc_0_5_ARID => twiddle_rsc_0_5_ARID,
      twiddle_rsc_0_5_BREADY => twiddle_rsc_0_5_BREADY,
      twiddle_rsc_0_5_BVALID => twiddle_rsc_0_5_BVALID,
      twiddle_rsc_0_5_BUSER => twiddle_rsc_0_5_BUSER,
      twiddle_rsc_0_5_BRESP => peaseNTT_core_inst_twiddle_rsc_0_5_BRESP,
      twiddle_rsc_0_5_BID => twiddle_rsc_0_5_BID,
      twiddle_rsc_0_5_WREADY => twiddle_rsc_0_5_WREADY,
      twiddle_rsc_0_5_WVALID => twiddle_rsc_0_5_WVALID,
      twiddle_rsc_0_5_WUSER => twiddle_rsc_0_5_WUSER,
      twiddle_rsc_0_5_WLAST => twiddle_rsc_0_5_WLAST,
      twiddle_rsc_0_5_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_5_WSTRB,
      twiddle_rsc_0_5_WDATA => peaseNTT_core_inst_twiddle_rsc_0_5_WDATA,
      twiddle_rsc_0_5_AWREADY => twiddle_rsc_0_5_AWREADY,
      twiddle_rsc_0_5_AWVALID => twiddle_rsc_0_5_AWVALID,
      twiddle_rsc_0_5_AWUSER => twiddle_rsc_0_5_AWUSER,
      twiddle_rsc_0_5_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_5_AWREGION,
      twiddle_rsc_0_5_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_5_AWQOS,
      twiddle_rsc_0_5_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_5_AWPROT,
      twiddle_rsc_0_5_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_5_AWCACHE,
      twiddle_rsc_0_5_AWLOCK => twiddle_rsc_0_5_AWLOCK,
      twiddle_rsc_0_5_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_5_AWBURST,
      twiddle_rsc_0_5_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_5_AWSIZE,
      twiddle_rsc_0_5_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_5_AWLEN,
      twiddle_rsc_0_5_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_5_AWADDR,
      twiddle_rsc_0_5_AWID => twiddle_rsc_0_5_AWID,
      twiddle_rsc_triosy_0_5_lz => twiddle_rsc_triosy_0_5_lz,
      twiddle_rsc_0_6_s_tdone => twiddle_rsc_0_6_s_tdone,
      twiddle_rsc_0_6_tr_write_done => twiddle_rsc_0_6_tr_write_done,
      twiddle_rsc_0_6_RREADY => twiddle_rsc_0_6_RREADY,
      twiddle_rsc_0_6_RVALID => twiddle_rsc_0_6_RVALID,
      twiddle_rsc_0_6_RUSER => twiddle_rsc_0_6_RUSER,
      twiddle_rsc_0_6_RLAST => twiddle_rsc_0_6_RLAST,
      twiddle_rsc_0_6_RRESP => peaseNTT_core_inst_twiddle_rsc_0_6_RRESP,
      twiddle_rsc_0_6_RDATA => peaseNTT_core_inst_twiddle_rsc_0_6_RDATA,
      twiddle_rsc_0_6_RID => twiddle_rsc_0_6_RID,
      twiddle_rsc_0_6_ARREADY => twiddle_rsc_0_6_ARREADY,
      twiddle_rsc_0_6_ARVALID => twiddle_rsc_0_6_ARVALID,
      twiddle_rsc_0_6_ARUSER => twiddle_rsc_0_6_ARUSER,
      twiddle_rsc_0_6_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_6_ARREGION,
      twiddle_rsc_0_6_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_6_ARQOS,
      twiddle_rsc_0_6_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_6_ARPROT,
      twiddle_rsc_0_6_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_6_ARCACHE,
      twiddle_rsc_0_6_ARLOCK => twiddle_rsc_0_6_ARLOCK,
      twiddle_rsc_0_6_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_6_ARBURST,
      twiddle_rsc_0_6_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_6_ARSIZE,
      twiddle_rsc_0_6_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_6_ARLEN,
      twiddle_rsc_0_6_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_6_ARADDR,
      twiddle_rsc_0_6_ARID => twiddle_rsc_0_6_ARID,
      twiddle_rsc_0_6_BREADY => twiddle_rsc_0_6_BREADY,
      twiddle_rsc_0_6_BVALID => twiddle_rsc_0_6_BVALID,
      twiddle_rsc_0_6_BUSER => twiddle_rsc_0_6_BUSER,
      twiddle_rsc_0_6_BRESP => peaseNTT_core_inst_twiddle_rsc_0_6_BRESP,
      twiddle_rsc_0_6_BID => twiddle_rsc_0_6_BID,
      twiddle_rsc_0_6_WREADY => twiddle_rsc_0_6_WREADY,
      twiddle_rsc_0_6_WVALID => twiddle_rsc_0_6_WVALID,
      twiddle_rsc_0_6_WUSER => twiddle_rsc_0_6_WUSER,
      twiddle_rsc_0_6_WLAST => twiddle_rsc_0_6_WLAST,
      twiddle_rsc_0_6_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_6_WSTRB,
      twiddle_rsc_0_6_WDATA => peaseNTT_core_inst_twiddle_rsc_0_6_WDATA,
      twiddle_rsc_0_6_AWREADY => twiddle_rsc_0_6_AWREADY,
      twiddle_rsc_0_6_AWVALID => twiddle_rsc_0_6_AWVALID,
      twiddle_rsc_0_6_AWUSER => twiddle_rsc_0_6_AWUSER,
      twiddle_rsc_0_6_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_6_AWREGION,
      twiddle_rsc_0_6_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_6_AWQOS,
      twiddle_rsc_0_6_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_6_AWPROT,
      twiddle_rsc_0_6_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_6_AWCACHE,
      twiddle_rsc_0_6_AWLOCK => twiddle_rsc_0_6_AWLOCK,
      twiddle_rsc_0_6_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_6_AWBURST,
      twiddle_rsc_0_6_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_6_AWSIZE,
      twiddle_rsc_0_6_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_6_AWLEN,
      twiddle_rsc_0_6_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_6_AWADDR,
      twiddle_rsc_0_6_AWID => twiddle_rsc_0_6_AWID,
      twiddle_rsc_triosy_0_6_lz => twiddle_rsc_triosy_0_6_lz,
      twiddle_rsc_0_7_s_tdone => twiddle_rsc_0_7_s_tdone,
      twiddle_rsc_0_7_tr_write_done => twiddle_rsc_0_7_tr_write_done,
      twiddle_rsc_0_7_RREADY => twiddle_rsc_0_7_RREADY,
      twiddle_rsc_0_7_RVALID => twiddle_rsc_0_7_RVALID,
      twiddle_rsc_0_7_RUSER => twiddle_rsc_0_7_RUSER,
      twiddle_rsc_0_7_RLAST => twiddle_rsc_0_7_RLAST,
      twiddle_rsc_0_7_RRESP => peaseNTT_core_inst_twiddle_rsc_0_7_RRESP,
      twiddle_rsc_0_7_RDATA => peaseNTT_core_inst_twiddle_rsc_0_7_RDATA,
      twiddle_rsc_0_7_RID => twiddle_rsc_0_7_RID,
      twiddle_rsc_0_7_ARREADY => twiddle_rsc_0_7_ARREADY,
      twiddle_rsc_0_7_ARVALID => twiddle_rsc_0_7_ARVALID,
      twiddle_rsc_0_7_ARUSER => twiddle_rsc_0_7_ARUSER,
      twiddle_rsc_0_7_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_7_ARREGION,
      twiddle_rsc_0_7_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_7_ARQOS,
      twiddle_rsc_0_7_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_7_ARPROT,
      twiddle_rsc_0_7_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_7_ARCACHE,
      twiddle_rsc_0_7_ARLOCK => twiddle_rsc_0_7_ARLOCK,
      twiddle_rsc_0_7_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_7_ARBURST,
      twiddle_rsc_0_7_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_7_ARSIZE,
      twiddle_rsc_0_7_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_7_ARLEN,
      twiddle_rsc_0_7_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_7_ARADDR,
      twiddle_rsc_0_7_ARID => twiddle_rsc_0_7_ARID,
      twiddle_rsc_0_7_BREADY => twiddle_rsc_0_7_BREADY,
      twiddle_rsc_0_7_BVALID => twiddle_rsc_0_7_BVALID,
      twiddle_rsc_0_7_BUSER => twiddle_rsc_0_7_BUSER,
      twiddle_rsc_0_7_BRESP => peaseNTT_core_inst_twiddle_rsc_0_7_BRESP,
      twiddle_rsc_0_7_BID => twiddle_rsc_0_7_BID,
      twiddle_rsc_0_7_WREADY => twiddle_rsc_0_7_WREADY,
      twiddle_rsc_0_7_WVALID => twiddle_rsc_0_7_WVALID,
      twiddle_rsc_0_7_WUSER => twiddle_rsc_0_7_WUSER,
      twiddle_rsc_0_7_WLAST => twiddle_rsc_0_7_WLAST,
      twiddle_rsc_0_7_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_7_WSTRB,
      twiddle_rsc_0_7_WDATA => peaseNTT_core_inst_twiddle_rsc_0_7_WDATA,
      twiddle_rsc_0_7_AWREADY => twiddle_rsc_0_7_AWREADY,
      twiddle_rsc_0_7_AWVALID => twiddle_rsc_0_7_AWVALID,
      twiddle_rsc_0_7_AWUSER => twiddle_rsc_0_7_AWUSER,
      twiddle_rsc_0_7_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_7_AWREGION,
      twiddle_rsc_0_7_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_7_AWQOS,
      twiddle_rsc_0_7_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_7_AWPROT,
      twiddle_rsc_0_7_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_7_AWCACHE,
      twiddle_rsc_0_7_AWLOCK => twiddle_rsc_0_7_AWLOCK,
      twiddle_rsc_0_7_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_7_AWBURST,
      twiddle_rsc_0_7_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_7_AWSIZE,
      twiddle_rsc_0_7_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_7_AWLEN,
      twiddle_rsc_0_7_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_7_AWADDR,
      twiddle_rsc_0_7_AWID => twiddle_rsc_0_7_AWID,
      twiddle_rsc_triosy_0_7_lz => twiddle_rsc_triosy_0_7_lz,
      twiddle_rsc_0_8_s_tdone => twiddle_rsc_0_8_s_tdone,
      twiddle_rsc_0_8_tr_write_done => twiddle_rsc_0_8_tr_write_done,
      twiddle_rsc_0_8_RREADY => twiddle_rsc_0_8_RREADY,
      twiddle_rsc_0_8_RVALID => twiddle_rsc_0_8_RVALID,
      twiddle_rsc_0_8_RUSER => twiddle_rsc_0_8_RUSER,
      twiddle_rsc_0_8_RLAST => twiddle_rsc_0_8_RLAST,
      twiddle_rsc_0_8_RRESP => peaseNTT_core_inst_twiddle_rsc_0_8_RRESP,
      twiddle_rsc_0_8_RDATA => peaseNTT_core_inst_twiddle_rsc_0_8_RDATA,
      twiddle_rsc_0_8_RID => twiddle_rsc_0_8_RID,
      twiddle_rsc_0_8_ARREADY => twiddle_rsc_0_8_ARREADY,
      twiddle_rsc_0_8_ARVALID => twiddle_rsc_0_8_ARVALID,
      twiddle_rsc_0_8_ARUSER => twiddle_rsc_0_8_ARUSER,
      twiddle_rsc_0_8_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_8_ARREGION,
      twiddle_rsc_0_8_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_8_ARQOS,
      twiddle_rsc_0_8_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_8_ARPROT,
      twiddle_rsc_0_8_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_8_ARCACHE,
      twiddle_rsc_0_8_ARLOCK => twiddle_rsc_0_8_ARLOCK,
      twiddle_rsc_0_8_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_8_ARBURST,
      twiddle_rsc_0_8_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_8_ARSIZE,
      twiddle_rsc_0_8_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_8_ARLEN,
      twiddle_rsc_0_8_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_8_ARADDR,
      twiddle_rsc_0_8_ARID => twiddle_rsc_0_8_ARID,
      twiddle_rsc_0_8_BREADY => twiddle_rsc_0_8_BREADY,
      twiddle_rsc_0_8_BVALID => twiddle_rsc_0_8_BVALID,
      twiddle_rsc_0_8_BUSER => twiddle_rsc_0_8_BUSER,
      twiddle_rsc_0_8_BRESP => peaseNTT_core_inst_twiddle_rsc_0_8_BRESP,
      twiddle_rsc_0_8_BID => twiddle_rsc_0_8_BID,
      twiddle_rsc_0_8_WREADY => twiddle_rsc_0_8_WREADY,
      twiddle_rsc_0_8_WVALID => twiddle_rsc_0_8_WVALID,
      twiddle_rsc_0_8_WUSER => twiddle_rsc_0_8_WUSER,
      twiddle_rsc_0_8_WLAST => twiddle_rsc_0_8_WLAST,
      twiddle_rsc_0_8_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_8_WSTRB,
      twiddle_rsc_0_8_WDATA => peaseNTT_core_inst_twiddle_rsc_0_8_WDATA,
      twiddle_rsc_0_8_AWREADY => twiddle_rsc_0_8_AWREADY,
      twiddle_rsc_0_8_AWVALID => twiddle_rsc_0_8_AWVALID,
      twiddle_rsc_0_8_AWUSER => twiddle_rsc_0_8_AWUSER,
      twiddle_rsc_0_8_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_8_AWREGION,
      twiddle_rsc_0_8_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_8_AWQOS,
      twiddle_rsc_0_8_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_8_AWPROT,
      twiddle_rsc_0_8_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_8_AWCACHE,
      twiddle_rsc_0_8_AWLOCK => twiddle_rsc_0_8_AWLOCK,
      twiddle_rsc_0_8_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_8_AWBURST,
      twiddle_rsc_0_8_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_8_AWSIZE,
      twiddle_rsc_0_8_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_8_AWLEN,
      twiddle_rsc_0_8_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_8_AWADDR,
      twiddle_rsc_0_8_AWID => twiddle_rsc_0_8_AWID,
      twiddle_rsc_triosy_0_8_lz => twiddle_rsc_triosy_0_8_lz,
      twiddle_rsc_0_9_s_tdone => twiddle_rsc_0_9_s_tdone,
      twiddle_rsc_0_9_tr_write_done => twiddle_rsc_0_9_tr_write_done,
      twiddle_rsc_0_9_RREADY => twiddle_rsc_0_9_RREADY,
      twiddle_rsc_0_9_RVALID => twiddle_rsc_0_9_RVALID,
      twiddle_rsc_0_9_RUSER => twiddle_rsc_0_9_RUSER,
      twiddle_rsc_0_9_RLAST => twiddle_rsc_0_9_RLAST,
      twiddle_rsc_0_9_RRESP => peaseNTT_core_inst_twiddle_rsc_0_9_RRESP,
      twiddle_rsc_0_9_RDATA => peaseNTT_core_inst_twiddle_rsc_0_9_RDATA,
      twiddle_rsc_0_9_RID => twiddle_rsc_0_9_RID,
      twiddle_rsc_0_9_ARREADY => twiddle_rsc_0_9_ARREADY,
      twiddle_rsc_0_9_ARVALID => twiddle_rsc_0_9_ARVALID,
      twiddle_rsc_0_9_ARUSER => twiddle_rsc_0_9_ARUSER,
      twiddle_rsc_0_9_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_9_ARREGION,
      twiddle_rsc_0_9_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_9_ARQOS,
      twiddle_rsc_0_9_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_9_ARPROT,
      twiddle_rsc_0_9_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_9_ARCACHE,
      twiddle_rsc_0_9_ARLOCK => twiddle_rsc_0_9_ARLOCK,
      twiddle_rsc_0_9_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_9_ARBURST,
      twiddle_rsc_0_9_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_9_ARSIZE,
      twiddle_rsc_0_9_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_9_ARLEN,
      twiddle_rsc_0_9_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_9_ARADDR,
      twiddle_rsc_0_9_ARID => twiddle_rsc_0_9_ARID,
      twiddle_rsc_0_9_BREADY => twiddle_rsc_0_9_BREADY,
      twiddle_rsc_0_9_BVALID => twiddle_rsc_0_9_BVALID,
      twiddle_rsc_0_9_BUSER => twiddle_rsc_0_9_BUSER,
      twiddle_rsc_0_9_BRESP => peaseNTT_core_inst_twiddle_rsc_0_9_BRESP,
      twiddle_rsc_0_9_BID => twiddle_rsc_0_9_BID,
      twiddle_rsc_0_9_WREADY => twiddle_rsc_0_9_WREADY,
      twiddle_rsc_0_9_WVALID => twiddle_rsc_0_9_WVALID,
      twiddle_rsc_0_9_WUSER => twiddle_rsc_0_9_WUSER,
      twiddle_rsc_0_9_WLAST => twiddle_rsc_0_9_WLAST,
      twiddle_rsc_0_9_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_9_WSTRB,
      twiddle_rsc_0_9_WDATA => peaseNTT_core_inst_twiddle_rsc_0_9_WDATA,
      twiddle_rsc_0_9_AWREADY => twiddle_rsc_0_9_AWREADY,
      twiddle_rsc_0_9_AWVALID => twiddle_rsc_0_9_AWVALID,
      twiddle_rsc_0_9_AWUSER => twiddle_rsc_0_9_AWUSER,
      twiddle_rsc_0_9_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_9_AWREGION,
      twiddle_rsc_0_9_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_9_AWQOS,
      twiddle_rsc_0_9_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_9_AWPROT,
      twiddle_rsc_0_9_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_9_AWCACHE,
      twiddle_rsc_0_9_AWLOCK => twiddle_rsc_0_9_AWLOCK,
      twiddle_rsc_0_9_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_9_AWBURST,
      twiddle_rsc_0_9_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_9_AWSIZE,
      twiddle_rsc_0_9_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_9_AWLEN,
      twiddle_rsc_0_9_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_9_AWADDR,
      twiddle_rsc_0_9_AWID => twiddle_rsc_0_9_AWID,
      twiddle_rsc_triosy_0_9_lz => twiddle_rsc_triosy_0_9_lz,
      twiddle_rsc_0_10_s_tdone => twiddle_rsc_0_10_s_tdone,
      twiddle_rsc_0_10_tr_write_done => twiddle_rsc_0_10_tr_write_done,
      twiddle_rsc_0_10_RREADY => twiddle_rsc_0_10_RREADY,
      twiddle_rsc_0_10_RVALID => twiddle_rsc_0_10_RVALID,
      twiddle_rsc_0_10_RUSER => twiddle_rsc_0_10_RUSER,
      twiddle_rsc_0_10_RLAST => twiddle_rsc_0_10_RLAST,
      twiddle_rsc_0_10_RRESP => peaseNTT_core_inst_twiddle_rsc_0_10_RRESP,
      twiddle_rsc_0_10_RDATA => peaseNTT_core_inst_twiddle_rsc_0_10_RDATA,
      twiddle_rsc_0_10_RID => twiddle_rsc_0_10_RID,
      twiddle_rsc_0_10_ARREADY => twiddle_rsc_0_10_ARREADY,
      twiddle_rsc_0_10_ARVALID => twiddle_rsc_0_10_ARVALID,
      twiddle_rsc_0_10_ARUSER => twiddle_rsc_0_10_ARUSER,
      twiddle_rsc_0_10_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_10_ARREGION,
      twiddle_rsc_0_10_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_10_ARQOS,
      twiddle_rsc_0_10_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_10_ARPROT,
      twiddle_rsc_0_10_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_10_ARCACHE,
      twiddle_rsc_0_10_ARLOCK => twiddle_rsc_0_10_ARLOCK,
      twiddle_rsc_0_10_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_10_ARBURST,
      twiddle_rsc_0_10_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_10_ARSIZE,
      twiddle_rsc_0_10_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_10_ARLEN,
      twiddle_rsc_0_10_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_10_ARADDR,
      twiddle_rsc_0_10_ARID => twiddle_rsc_0_10_ARID,
      twiddle_rsc_0_10_BREADY => twiddle_rsc_0_10_BREADY,
      twiddle_rsc_0_10_BVALID => twiddle_rsc_0_10_BVALID,
      twiddle_rsc_0_10_BUSER => twiddle_rsc_0_10_BUSER,
      twiddle_rsc_0_10_BRESP => peaseNTT_core_inst_twiddle_rsc_0_10_BRESP,
      twiddle_rsc_0_10_BID => twiddle_rsc_0_10_BID,
      twiddle_rsc_0_10_WREADY => twiddle_rsc_0_10_WREADY,
      twiddle_rsc_0_10_WVALID => twiddle_rsc_0_10_WVALID,
      twiddle_rsc_0_10_WUSER => twiddle_rsc_0_10_WUSER,
      twiddle_rsc_0_10_WLAST => twiddle_rsc_0_10_WLAST,
      twiddle_rsc_0_10_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_10_WSTRB,
      twiddle_rsc_0_10_WDATA => peaseNTT_core_inst_twiddle_rsc_0_10_WDATA,
      twiddle_rsc_0_10_AWREADY => twiddle_rsc_0_10_AWREADY,
      twiddle_rsc_0_10_AWVALID => twiddle_rsc_0_10_AWVALID,
      twiddle_rsc_0_10_AWUSER => twiddle_rsc_0_10_AWUSER,
      twiddle_rsc_0_10_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_10_AWREGION,
      twiddle_rsc_0_10_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_10_AWQOS,
      twiddle_rsc_0_10_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_10_AWPROT,
      twiddle_rsc_0_10_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_10_AWCACHE,
      twiddle_rsc_0_10_AWLOCK => twiddle_rsc_0_10_AWLOCK,
      twiddle_rsc_0_10_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_10_AWBURST,
      twiddle_rsc_0_10_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_10_AWSIZE,
      twiddle_rsc_0_10_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_10_AWLEN,
      twiddle_rsc_0_10_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_10_AWADDR,
      twiddle_rsc_0_10_AWID => twiddle_rsc_0_10_AWID,
      twiddle_rsc_triosy_0_10_lz => twiddle_rsc_triosy_0_10_lz,
      twiddle_rsc_0_11_s_tdone => twiddle_rsc_0_11_s_tdone,
      twiddle_rsc_0_11_tr_write_done => twiddle_rsc_0_11_tr_write_done,
      twiddle_rsc_0_11_RREADY => twiddle_rsc_0_11_RREADY,
      twiddle_rsc_0_11_RVALID => twiddle_rsc_0_11_RVALID,
      twiddle_rsc_0_11_RUSER => twiddle_rsc_0_11_RUSER,
      twiddle_rsc_0_11_RLAST => twiddle_rsc_0_11_RLAST,
      twiddle_rsc_0_11_RRESP => peaseNTT_core_inst_twiddle_rsc_0_11_RRESP,
      twiddle_rsc_0_11_RDATA => peaseNTT_core_inst_twiddle_rsc_0_11_RDATA,
      twiddle_rsc_0_11_RID => twiddle_rsc_0_11_RID,
      twiddle_rsc_0_11_ARREADY => twiddle_rsc_0_11_ARREADY,
      twiddle_rsc_0_11_ARVALID => twiddle_rsc_0_11_ARVALID,
      twiddle_rsc_0_11_ARUSER => twiddle_rsc_0_11_ARUSER,
      twiddle_rsc_0_11_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_11_ARREGION,
      twiddle_rsc_0_11_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_11_ARQOS,
      twiddle_rsc_0_11_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_11_ARPROT,
      twiddle_rsc_0_11_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_11_ARCACHE,
      twiddle_rsc_0_11_ARLOCK => twiddle_rsc_0_11_ARLOCK,
      twiddle_rsc_0_11_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_11_ARBURST,
      twiddle_rsc_0_11_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_11_ARSIZE,
      twiddle_rsc_0_11_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_11_ARLEN,
      twiddle_rsc_0_11_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_11_ARADDR,
      twiddle_rsc_0_11_ARID => twiddle_rsc_0_11_ARID,
      twiddle_rsc_0_11_BREADY => twiddle_rsc_0_11_BREADY,
      twiddle_rsc_0_11_BVALID => twiddle_rsc_0_11_BVALID,
      twiddle_rsc_0_11_BUSER => twiddle_rsc_0_11_BUSER,
      twiddle_rsc_0_11_BRESP => peaseNTT_core_inst_twiddle_rsc_0_11_BRESP,
      twiddle_rsc_0_11_BID => twiddle_rsc_0_11_BID,
      twiddle_rsc_0_11_WREADY => twiddle_rsc_0_11_WREADY,
      twiddle_rsc_0_11_WVALID => twiddle_rsc_0_11_WVALID,
      twiddle_rsc_0_11_WUSER => twiddle_rsc_0_11_WUSER,
      twiddle_rsc_0_11_WLAST => twiddle_rsc_0_11_WLAST,
      twiddle_rsc_0_11_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_11_WSTRB,
      twiddle_rsc_0_11_WDATA => peaseNTT_core_inst_twiddle_rsc_0_11_WDATA,
      twiddle_rsc_0_11_AWREADY => twiddle_rsc_0_11_AWREADY,
      twiddle_rsc_0_11_AWVALID => twiddle_rsc_0_11_AWVALID,
      twiddle_rsc_0_11_AWUSER => twiddle_rsc_0_11_AWUSER,
      twiddle_rsc_0_11_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_11_AWREGION,
      twiddle_rsc_0_11_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_11_AWQOS,
      twiddle_rsc_0_11_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_11_AWPROT,
      twiddle_rsc_0_11_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_11_AWCACHE,
      twiddle_rsc_0_11_AWLOCK => twiddle_rsc_0_11_AWLOCK,
      twiddle_rsc_0_11_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_11_AWBURST,
      twiddle_rsc_0_11_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_11_AWSIZE,
      twiddle_rsc_0_11_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_11_AWLEN,
      twiddle_rsc_0_11_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_11_AWADDR,
      twiddle_rsc_0_11_AWID => twiddle_rsc_0_11_AWID,
      twiddle_rsc_triosy_0_11_lz => twiddle_rsc_triosy_0_11_lz,
      twiddle_rsc_0_12_s_tdone => twiddle_rsc_0_12_s_tdone,
      twiddle_rsc_0_12_tr_write_done => twiddle_rsc_0_12_tr_write_done,
      twiddle_rsc_0_12_RREADY => twiddle_rsc_0_12_RREADY,
      twiddle_rsc_0_12_RVALID => twiddle_rsc_0_12_RVALID,
      twiddle_rsc_0_12_RUSER => twiddle_rsc_0_12_RUSER,
      twiddle_rsc_0_12_RLAST => twiddle_rsc_0_12_RLAST,
      twiddle_rsc_0_12_RRESP => peaseNTT_core_inst_twiddle_rsc_0_12_RRESP,
      twiddle_rsc_0_12_RDATA => peaseNTT_core_inst_twiddle_rsc_0_12_RDATA,
      twiddle_rsc_0_12_RID => twiddle_rsc_0_12_RID,
      twiddle_rsc_0_12_ARREADY => twiddle_rsc_0_12_ARREADY,
      twiddle_rsc_0_12_ARVALID => twiddle_rsc_0_12_ARVALID,
      twiddle_rsc_0_12_ARUSER => twiddle_rsc_0_12_ARUSER,
      twiddle_rsc_0_12_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_12_ARREGION,
      twiddle_rsc_0_12_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_12_ARQOS,
      twiddle_rsc_0_12_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_12_ARPROT,
      twiddle_rsc_0_12_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_12_ARCACHE,
      twiddle_rsc_0_12_ARLOCK => twiddle_rsc_0_12_ARLOCK,
      twiddle_rsc_0_12_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_12_ARBURST,
      twiddle_rsc_0_12_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_12_ARSIZE,
      twiddle_rsc_0_12_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_12_ARLEN,
      twiddle_rsc_0_12_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_12_ARADDR,
      twiddle_rsc_0_12_ARID => twiddle_rsc_0_12_ARID,
      twiddle_rsc_0_12_BREADY => twiddle_rsc_0_12_BREADY,
      twiddle_rsc_0_12_BVALID => twiddle_rsc_0_12_BVALID,
      twiddle_rsc_0_12_BUSER => twiddle_rsc_0_12_BUSER,
      twiddle_rsc_0_12_BRESP => peaseNTT_core_inst_twiddle_rsc_0_12_BRESP,
      twiddle_rsc_0_12_BID => twiddle_rsc_0_12_BID,
      twiddle_rsc_0_12_WREADY => twiddle_rsc_0_12_WREADY,
      twiddle_rsc_0_12_WVALID => twiddle_rsc_0_12_WVALID,
      twiddle_rsc_0_12_WUSER => twiddle_rsc_0_12_WUSER,
      twiddle_rsc_0_12_WLAST => twiddle_rsc_0_12_WLAST,
      twiddle_rsc_0_12_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_12_WSTRB,
      twiddle_rsc_0_12_WDATA => peaseNTT_core_inst_twiddle_rsc_0_12_WDATA,
      twiddle_rsc_0_12_AWREADY => twiddle_rsc_0_12_AWREADY,
      twiddle_rsc_0_12_AWVALID => twiddle_rsc_0_12_AWVALID,
      twiddle_rsc_0_12_AWUSER => twiddle_rsc_0_12_AWUSER,
      twiddle_rsc_0_12_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_12_AWREGION,
      twiddle_rsc_0_12_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_12_AWQOS,
      twiddle_rsc_0_12_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_12_AWPROT,
      twiddle_rsc_0_12_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_12_AWCACHE,
      twiddle_rsc_0_12_AWLOCK => twiddle_rsc_0_12_AWLOCK,
      twiddle_rsc_0_12_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_12_AWBURST,
      twiddle_rsc_0_12_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_12_AWSIZE,
      twiddle_rsc_0_12_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_12_AWLEN,
      twiddle_rsc_0_12_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_12_AWADDR,
      twiddle_rsc_0_12_AWID => twiddle_rsc_0_12_AWID,
      twiddle_rsc_triosy_0_12_lz => twiddle_rsc_triosy_0_12_lz,
      twiddle_rsc_0_13_s_tdone => twiddle_rsc_0_13_s_tdone,
      twiddle_rsc_0_13_tr_write_done => twiddle_rsc_0_13_tr_write_done,
      twiddle_rsc_0_13_RREADY => twiddle_rsc_0_13_RREADY,
      twiddle_rsc_0_13_RVALID => twiddle_rsc_0_13_RVALID,
      twiddle_rsc_0_13_RUSER => twiddle_rsc_0_13_RUSER,
      twiddle_rsc_0_13_RLAST => twiddle_rsc_0_13_RLAST,
      twiddle_rsc_0_13_RRESP => peaseNTT_core_inst_twiddle_rsc_0_13_RRESP,
      twiddle_rsc_0_13_RDATA => peaseNTT_core_inst_twiddle_rsc_0_13_RDATA,
      twiddle_rsc_0_13_RID => twiddle_rsc_0_13_RID,
      twiddle_rsc_0_13_ARREADY => twiddle_rsc_0_13_ARREADY,
      twiddle_rsc_0_13_ARVALID => twiddle_rsc_0_13_ARVALID,
      twiddle_rsc_0_13_ARUSER => twiddle_rsc_0_13_ARUSER,
      twiddle_rsc_0_13_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_13_ARREGION,
      twiddle_rsc_0_13_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_13_ARQOS,
      twiddle_rsc_0_13_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_13_ARPROT,
      twiddle_rsc_0_13_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_13_ARCACHE,
      twiddle_rsc_0_13_ARLOCK => twiddle_rsc_0_13_ARLOCK,
      twiddle_rsc_0_13_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_13_ARBURST,
      twiddle_rsc_0_13_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_13_ARSIZE,
      twiddle_rsc_0_13_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_13_ARLEN,
      twiddle_rsc_0_13_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_13_ARADDR,
      twiddle_rsc_0_13_ARID => twiddle_rsc_0_13_ARID,
      twiddle_rsc_0_13_BREADY => twiddle_rsc_0_13_BREADY,
      twiddle_rsc_0_13_BVALID => twiddle_rsc_0_13_BVALID,
      twiddle_rsc_0_13_BUSER => twiddle_rsc_0_13_BUSER,
      twiddle_rsc_0_13_BRESP => peaseNTT_core_inst_twiddle_rsc_0_13_BRESP,
      twiddle_rsc_0_13_BID => twiddle_rsc_0_13_BID,
      twiddle_rsc_0_13_WREADY => twiddle_rsc_0_13_WREADY,
      twiddle_rsc_0_13_WVALID => twiddle_rsc_0_13_WVALID,
      twiddle_rsc_0_13_WUSER => twiddle_rsc_0_13_WUSER,
      twiddle_rsc_0_13_WLAST => twiddle_rsc_0_13_WLAST,
      twiddle_rsc_0_13_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_13_WSTRB,
      twiddle_rsc_0_13_WDATA => peaseNTT_core_inst_twiddle_rsc_0_13_WDATA,
      twiddle_rsc_0_13_AWREADY => twiddle_rsc_0_13_AWREADY,
      twiddle_rsc_0_13_AWVALID => twiddle_rsc_0_13_AWVALID,
      twiddle_rsc_0_13_AWUSER => twiddle_rsc_0_13_AWUSER,
      twiddle_rsc_0_13_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_13_AWREGION,
      twiddle_rsc_0_13_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_13_AWQOS,
      twiddle_rsc_0_13_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_13_AWPROT,
      twiddle_rsc_0_13_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_13_AWCACHE,
      twiddle_rsc_0_13_AWLOCK => twiddle_rsc_0_13_AWLOCK,
      twiddle_rsc_0_13_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_13_AWBURST,
      twiddle_rsc_0_13_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_13_AWSIZE,
      twiddle_rsc_0_13_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_13_AWLEN,
      twiddle_rsc_0_13_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_13_AWADDR,
      twiddle_rsc_0_13_AWID => twiddle_rsc_0_13_AWID,
      twiddle_rsc_triosy_0_13_lz => twiddle_rsc_triosy_0_13_lz,
      twiddle_rsc_0_14_s_tdone => twiddle_rsc_0_14_s_tdone,
      twiddle_rsc_0_14_tr_write_done => twiddle_rsc_0_14_tr_write_done,
      twiddle_rsc_0_14_RREADY => twiddle_rsc_0_14_RREADY,
      twiddle_rsc_0_14_RVALID => twiddle_rsc_0_14_RVALID,
      twiddle_rsc_0_14_RUSER => twiddle_rsc_0_14_RUSER,
      twiddle_rsc_0_14_RLAST => twiddle_rsc_0_14_RLAST,
      twiddle_rsc_0_14_RRESP => peaseNTT_core_inst_twiddle_rsc_0_14_RRESP,
      twiddle_rsc_0_14_RDATA => peaseNTT_core_inst_twiddle_rsc_0_14_RDATA,
      twiddle_rsc_0_14_RID => twiddle_rsc_0_14_RID,
      twiddle_rsc_0_14_ARREADY => twiddle_rsc_0_14_ARREADY,
      twiddle_rsc_0_14_ARVALID => twiddle_rsc_0_14_ARVALID,
      twiddle_rsc_0_14_ARUSER => twiddle_rsc_0_14_ARUSER,
      twiddle_rsc_0_14_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_14_ARREGION,
      twiddle_rsc_0_14_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_14_ARQOS,
      twiddle_rsc_0_14_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_14_ARPROT,
      twiddle_rsc_0_14_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_14_ARCACHE,
      twiddle_rsc_0_14_ARLOCK => twiddle_rsc_0_14_ARLOCK,
      twiddle_rsc_0_14_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_14_ARBURST,
      twiddle_rsc_0_14_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_14_ARSIZE,
      twiddle_rsc_0_14_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_14_ARLEN,
      twiddle_rsc_0_14_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_14_ARADDR,
      twiddle_rsc_0_14_ARID => twiddle_rsc_0_14_ARID,
      twiddle_rsc_0_14_BREADY => twiddle_rsc_0_14_BREADY,
      twiddle_rsc_0_14_BVALID => twiddle_rsc_0_14_BVALID,
      twiddle_rsc_0_14_BUSER => twiddle_rsc_0_14_BUSER,
      twiddle_rsc_0_14_BRESP => peaseNTT_core_inst_twiddle_rsc_0_14_BRESP,
      twiddle_rsc_0_14_BID => twiddle_rsc_0_14_BID,
      twiddle_rsc_0_14_WREADY => twiddle_rsc_0_14_WREADY,
      twiddle_rsc_0_14_WVALID => twiddle_rsc_0_14_WVALID,
      twiddle_rsc_0_14_WUSER => twiddle_rsc_0_14_WUSER,
      twiddle_rsc_0_14_WLAST => twiddle_rsc_0_14_WLAST,
      twiddle_rsc_0_14_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_14_WSTRB,
      twiddle_rsc_0_14_WDATA => peaseNTT_core_inst_twiddle_rsc_0_14_WDATA,
      twiddle_rsc_0_14_AWREADY => twiddle_rsc_0_14_AWREADY,
      twiddle_rsc_0_14_AWVALID => twiddle_rsc_0_14_AWVALID,
      twiddle_rsc_0_14_AWUSER => twiddle_rsc_0_14_AWUSER,
      twiddle_rsc_0_14_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_14_AWREGION,
      twiddle_rsc_0_14_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_14_AWQOS,
      twiddle_rsc_0_14_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_14_AWPROT,
      twiddle_rsc_0_14_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_14_AWCACHE,
      twiddle_rsc_0_14_AWLOCK => twiddle_rsc_0_14_AWLOCK,
      twiddle_rsc_0_14_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_14_AWBURST,
      twiddle_rsc_0_14_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_14_AWSIZE,
      twiddle_rsc_0_14_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_14_AWLEN,
      twiddle_rsc_0_14_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_14_AWADDR,
      twiddle_rsc_0_14_AWID => twiddle_rsc_0_14_AWID,
      twiddle_rsc_triosy_0_14_lz => twiddle_rsc_triosy_0_14_lz,
      twiddle_rsc_0_15_s_tdone => twiddle_rsc_0_15_s_tdone,
      twiddle_rsc_0_15_tr_write_done => twiddle_rsc_0_15_tr_write_done,
      twiddle_rsc_0_15_RREADY => twiddle_rsc_0_15_RREADY,
      twiddle_rsc_0_15_RVALID => twiddle_rsc_0_15_RVALID,
      twiddle_rsc_0_15_RUSER => twiddle_rsc_0_15_RUSER,
      twiddle_rsc_0_15_RLAST => twiddle_rsc_0_15_RLAST,
      twiddle_rsc_0_15_RRESP => peaseNTT_core_inst_twiddle_rsc_0_15_RRESP,
      twiddle_rsc_0_15_RDATA => peaseNTT_core_inst_twiddle_rsc_0_15_RDATA,
      twiddle_rsc_0_15_RID => twiddle_rsc_0_15_RID,
      twiddle_rsc_0_15_ARREADY => twiddle_rsc_0_15_ARREADY,
      twiddle_rsc_0_15_ARVALID => twiddle_rsc_0_15_ARVALID,
      twiddle_rsc_0_15_ARUSER => twiddle_rsc_0_15_ARUSER,
      twiddle_rsc_0_15_ARREGION => peaseNTT_core_inst_twiddle_rsc_0_15_ARREGION,
      twiddle_rsc_0_15_ARQOS => peaseNTT_core_inst_twiddle_rsc_0_15_ARQOS,
      twiddle_rsc_0_15_ARPROT => peaseNTT_core_inst_twiddle_rsc_0_15_ARPROT,
      twiddle_rsc_0_15_ARCACHE => peaseNTT_core_inst_twiddle_rsc_0_15_ARCACHE,
      twiddle_rsc_0_15_ARLOCK => twiddle_rsc_0_15_ARLOCK,
      twiddle_rsc_0_15_ARBURST => peaseNTT_core_inst_twiddle_rsc_0_15_ARBURST,
      twiddle_rsc_0_15_ARSIZE => peaseNTT_core_inst_twiddle_rsc_0_15_ARSIZE,
      twiddle_rsc_0_15_ARLEN => peaseNTT_core_inst_twiddle_rsc_0_15_ARLEN,
      twiddle_rsc_0_15_ARADDR => peaseNTT_core_inst_twiddle_rsc_0_15_ARADDR,
      twiddle_rsc_0_15_ARID => twiddle_rsc_0_15_ARID,
      twiddle_rsc_0_15_BREADY => twiddle_rsc_0_15_BREADY,
      twiddle_rsc_0_15_BVALID => twiddle_rsc_0_15_BVALID,
      twiddle_rsc_0_15_BUSER => twiddle_rsc_0_15_BUSER,
      twiddle_rsc_0_15_BRESP => peaseNTT_core_inst_twiddle_rsc_0_15_BRESP,
      twiddle_rsc_0_15_BID => twiddle_rsc_0_15_BID,
      twiddle_rsc_0_15_WREADY => twiddle_rsc_0_15_WREADY,
      twiddle_rsc_0_15_WVALID => twiddle_rsc_0_15_WVALID,
      twiddle_rsc_0_15_WUSER => twiddle_rsc_0_15_WUSER,
      twiddle_rsc_0_15_WLAST => twiddle_rsc_0_15_WLAST,
      twiddle_rsc_0_15_WSTRB => peaseNTT_core_inst_twiddle_rsc_0_15_WSTRB,
      twiddle_rsc_0_15_WDATA => peaseNTT_core_inst_twiddle_rsc_0_15_WDATA,
      twiddle_rsc_0_15_AWREADY => twiddle_rsc_0_15_AWREADY,
      twiddle_rsc_0_15_AWVALID => twiddle_rsc_0_15_AWVALID,
      twiddle_rsc_0_15_AWUSER => twiddle_rsc_0_15_AWUSER,
      twiddle_rsc_0_15_AWREGION => peaseNTT_core_inst_twiddle_rsc_0_15_AWREGION,
      twiddle_rsc_0_15_AWQOS => peaseNTT_core_inst_twiddle_rsc_0_15_AWQOS,
      twiddle_rsc_0_15_AWPROT => peaseNTT_core_inst_twiddle_rsc_0_15_AWPROT,
      twiddle_rsc_0_15_AWCACHE => peaseNTT_core_inst_twiddle_rsc_0_15_AWCACHE,
      twiddle_rsc_0_15_AWLOCK => twiddle_rsc_0_15_AWLOCK,
      twiddle_rsc_0_15_AWBURST => peaseNTT_core_inst_twiddle_rsc_0_15_AWBURST,
      twiddle_rsc_0_15_AWSIZE => peaseNTT_core_inst_twiddle_rsc_0_15_AWSIZE,
      twiddle_rsc_0_15_AWLEN => peaseNTT_core_inst_twiddle_rsc_0_15_AWLEN,
      twiddle_rsc_0_15_AWADDR => peaseNTT_core_inst_twiddle_rsc_0_15_AWADDR,
      twiddle_rsc_0_15_AWID => twiddle_rsc_0_15_AWID,
      twiddle_rsc_triosy_0_15_lz => twiddle_rsc_triosy_0_15_lz,
      twiddle_h_rsc_0_0_s_tdone => twiddle_h_rsc_0_0_s_tdone,
      twiddle_h_rsc_0_0_tr_write_done => twiddle_h_rsc_0_0_tr_write_done,
      twiddle_h_rsc_0_0_RREADY => twiddle_h_rsc_0_0_RREADY,
      twiddle_h_rsc_0_0_RVALID => twiddle_h_rsc_0_0_RVALID,
      twiddle_h_rsc_0_0_RUSER => twiddle_h_rsc_0_0_RUSER,
      twiddle_h_rsc_0_0_RLAST => twiddle_h_rsc_0_0_RLAST,
      twiddle_h_rsc_0_0_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_0_RRESP,
      twiddle_h_rsc_0_0_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_0_RDATA,
      twiddle_h_rsc_0_0_RID => twiddle_h_rsc_0_0_RID,
      twiddle_h_rsc_0_0_ARREADY => twiddle_h_rsc_0_0_ARREADY,
      twiddle_h_rsc_0_0_ARVALID => twiddle_h_rsc_0_0_ARVALID,
      twiddle_h_rsc_0_0_ARUSER => twiddle_h_rsc_0_0_ARUSER,
      twiddle_h_rsc_0_0_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_0_ARREGION,
      twiddle_h_rsc_0_0_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_0_ARQOS,
      twiddle_h_rsc_0_0_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_0_ARPROT,
      twiddle_h_rsc_0_0_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_0_ARCACHE,
      twiddle_h_rsc_0_0_ARLOCK => twiddle_h_rsc_0_0_ARLOCK,
      twiddle_h_rsc_0_0_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_0_ARBURST,
      twiddle_h_rsc_0_0_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_0_ARSIZE,
      twiddle_h_rsc_0_0_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_0_ARLEN,
      twiddle_h_rsc_0_0_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_0_ARADDR,
      twiddle_h_rsc_0_0_ARID => twiddle_h_rsc_0_0_ARID,
      twiddle_h_rsc_0_0_BREADY => twiddle_h_rsc_0_0_BREADY,
      twiddle_h_rsc_0_0_BVALID => twiddle_h_rsc_0_0_BVALID,
      twiddle_h_rsc_0_0_BUSER => twiddle_h_rsc_0_0_BUSER,
      twiddle_h_rsc_0_0_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_0_BRESP,
      twiddle_h_rsc_0_0_BID => twiddle_h_rsc_0_0_BID,
      twiddle_h_rsc_0_0_WREADY => twiddle_h_rsc_0_0_WREADY,
      twiddle_h_rsc_0_0_WVALID => twiddle_h_rsc_0_0_WVALID,
      twiddle_h_rsc_0_0_WUSER => twiddle_h_rsc_0_0_WUSER,
      twiddle_h_rsc_0_0_WLAST => twiddle_h_rsc_0_0_WLAST,
      twiddle_h_rsc_0_0_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_0_WSTRB,
      twiddle_h_rsc_0_0_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_0_WDATA,
      twiddle_h_rsc_0_0_AWREADY => twiddle_h_rsc_0_0_AWREADY,
      twiddle_h_rsc_0_0_AWVALID => twiddle_h_rsc_0_0_AWVALID,
      twiddle_h_rsc_0_0_AWUSER => twiddle_h_rsc_0_0_AWUSER,
      twiddle_h_rsc_0_0_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_0_AWREGION,
      twiddle_h_rsc_0_0_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_0_AWQOS,
      twiddle_h_rsc_0_0_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_0_AWPROT,
      twiddle_h_rsc_0_0_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_0_AWCACHE,
      twiddle_h_rsc_0_0_AWLOCK => twiddle_h_rsc_0_0_AWLOCK,
      twiddle_h_rsc_0_0_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_0_AWBURST,
      twiddle_h_rsc_0_0_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_0_AWSIZE,
      twiddle_h_rsc_0_0_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_0_AWLEN,
      twiddle_h_rsc_0_0_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_0_AWADDR,
      twiddle_h_rsc_0_0_AWID => twiddle_h_rsc_0_0_AWID,
      twiddle_h_rsc_triosy_0_0_lz => twiddle_h_rsc_triosy_0_0_lz,
      twiddle_h_rsc_0_1_s_tdone => twiddle_h_rsc_0_1_s_tdone,
      twiddle_h_rsc_0_1_tr_write_done => twiddle_h_rsc_0_1_tr_write_done,
      twiddle_h_rsc_0_1_RREADY => twiddle_h_rsc_0_1_RREADY,
      twiddle_h_rsc_0_1_RVALID => twiddle_h_rsc_0_1_RVALID,
      twiddle_h_rsc_0_1_RUSER => twiddle_h_rsc_0_1_RUSER,
      twiddle_h_rsc_0_1_RLAST => twiddle_h_rsc_0_1_RLAST,
      twiddle_h_rsc_0_1_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_1_RRESP,
      twiddle_h_rsc_0_1_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_1_RDATA,
      twiddle_h_rsc_0_1_RID => twiddle_h_rsc_0_1_RID,
      twiddle_h_rsc_0_1_ARREADY => twiddle_h_rsc_0_1_ARREADY,
      twiddle_h_rsc_0_1_ARVALID => twiddle_h_rsc_0_1_ARVALID,
      twiddle_h_rsc_0_1_ARUSER => twiddle_h_rsc_0_1_ARUSER,
      twiddle_h_rsc_0_1_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_1_ARREGION,
      twiddle_h_rsc_0_1_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_1_ARQOS,
      twiddle_h_rsc_0_1_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_1_ARPROT,
      twiddle_h_rsc_0_1_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_1_ARCACHE,
      twiddle_h_rsc_0_1_ARLOCK => twiddle_h_rsc_0_1_ARLOCK,
      twiddle_h_rsc_0_1_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_1_ARBURST,
      twiddle_h_rsc_0_1_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_1_ARSIZE,
      twiddle_h_rsc_0_1_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_1_ARLEN,
      twiddle_h_rsc_0_1_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_1_ARADDR,
      twiddle_h_rsc_0_1_ARID => twiddle_h_rsc_0_1_ARID,
      twiddle_h_rsc_0_1_BREADY => twiddle_h_rsc_0_1_BREADY,
      twiddle_h_rsc_0_1_BVALID => twiddle_h_rsc_0_1_BVALID,
      twiddle_h_rsc_0_1_BUSER => twiddle_h_rsc_0_1_BUSER,
      twiddle_h_rsc_0_1_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_1_BRESP,
      twiddle_h_rsc_0_1_BID => twiddle_h_rsc_0_1_BID,
      twiddle_h_rsc_0_1_WREADY => twiddle_h_rsc_0_1_WREADY,
      twiddle_h_rsc_0_1_WVALID => twiddle_h_rsc_0_1_WVALID,
      twiddle_h_rsc_0_1_WUSER => twiddle_h_rsc_0_1_WUSER,
      twiddle_h_rsc_0_1_WLAST => twiddle_h_rsc_0_1_WLAST,
      twiddle_h_rsc_0_1_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_1_WSTRB,
      twiddle_h_rsc_0_1_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_1_WDATA,
      twiddle_h_rsc_0_1_AWREADY => twiddle_h_rsc_0_1_AWREADY,
      twiddle_h_rsc_0_1_AWVALID => twiddle_h_rsc_0_1_AWVALID,
      twiddle_h_rsc_0_1_AWUSER => twiddle_h_rsc_0_1_AWUSER,
      twiddle_h_rsc_0_1_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_1_AWREGION,
      twiddle_h_rsc_0_1_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_1_AWQOS,
      twiddle_h_rsc_0_1_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_1_AWPROT,
      twiddle_h_rsc_0_1_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_1_AWCACHE,
      twiddle_h_rsc_0_1_AWLOCK => twiddle_h_rsc_0_1_AWLOCK,
      twiddle_h_rsc_0_1_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_1_AWBURST,
      twiddle_h_rsc_0_1_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_1_AWSIZE,
      twiddle_h_rsc_0_1_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_1_AWLEN,
      twiddle_h_rsc_0_1_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_1_AWADDR,
      twiddle_h_rsc_0_1_AWID => twiddle_h_rsc_0_1_AWID,
      twiddle_h_rsc_triosy_0_1_lz => twiddle_h_rsc_triosy_0_1_lz,
      twiddle_h_rsc_0_2_s_tdone => twiddle_h_rsc_0_2_s_tdone,
      twiddle_h_rsc_0_2_tr_write_done => twiddle_h_rsc_0_2_tr_write_done,
      twiddle_h_rsc_0_2_RREADY => twiddle_h_rsc_0_2_RREADY,
      twiddle_h_rsc_0_2_RVALID => twiddle_h_rsc_0_2_RVALID,
      twiddle_h_rsc_0_2_RUSER => twiddle_h_rsc_0_2_RUSER,
      twiddle_h_rsc_0_2_RLAST => twiddle_h_rsc_0_2_RLAST,
      twiddle_h_rsc_0_2_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_2_RRESP,
      twiddle_h_rsc_0_2_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_2_RDATA,
      twiddle_h_rsc_0_2_RID => twiddle_h_rsc_0_2_RID,
      twiddle_h_rsc_0_2_ARREADY => twiddle_h_rsc_0_2_ARREADY,
      twiddle_h_rsc_0_2_ARVALID => twiddle_h_rsc_0_2_ARVALID,
      twiddle_h_rsc_0_2_ARUSER => twiddle_h_rsc_0_2_ARUSER,
      twiddle_h_rsc_0_2_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_2_ARREGION,
      twiddle_h_rsc_0_2_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_2_ARQOS,
      twiddle_h_rsc_0_2_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_2_ARPROT,
      twiddle_h_rsc_0_2_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_2_ARCACHE,
      twiddle_h_rsc_0_2_ARLOCK => twiddle_h_rsc_0_2_ARLOCK,
      twiddle_h_rsc_0_2_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_2_ARBURST,
      twiddle_h_rsc_0_2_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_2_ARSIZE,
      twiddle_h_rsc_0_2_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_2_ARLEN,
      twiddle_h_rsc_0_2_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_2_ARADDR,
      twiddle_h_rsc_0_2_ARID => twiddle_h_rsc_0_2_ARID,
      twiddle_h_rsc_0_2_BREADY => twiddle_h_rsc_0_2_BREADY,
      twiddle_h_rsc_0_2_BVALID => twiddle_h_rsc_0_2_BVALID,
      twiddle_h_rsc_0_2_BUSER => twiddle_h_rsc_0_2_BUSER,
      twiddle_h_rsc_0_2_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_2_BRESP,
      twiddle_h_rsc_0_2_BID => twiddle_h_rsc_0_2_BID,
      twiddle_h_rsc_0_2_WREADY => twiddle_h_rsc_0_2_WREADY,
      twiddle_h_rsc_0_2_WVALID => twiddle_h_rsc_0_2_WVALID,
      twiddle_h_rsc_0_2_WUSER => twiddle_h_rsc_0_2_WUSER,
      twiddle_h_rsc_0_2_WLAST => twiddle_h_rsc_0_2_WLAST,
      twiddle_h_rsc_0_2_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_2_WSTRB,
      twiddle_h_rsc_0_2_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_2_WDATA,
      twiddle_h_rsc_0_2_AWREADY => twiddle_h_rsc_0_2_AWREADY,
      twiddle_h_rsc_0_2_AWVALID => twiddle_h_rsc_0_2_AWVALID,
      twiddle_h_rsc_0_2_AWUSER => twiddle_h_rsc_0_2_AWUSER,
      twiddle_h_rsc_0_2_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_2_AWREGION,
      twiddle_h_rsc_0_2_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_2_AWQOS,
      twiddle_h_rsc_0_2_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_2_AWPROT,
      twiddle_h_rsc_0_2_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_2_AWCACHE,
      twiddle_h_rsc_0_2_AWLOCK => twiddle_h_rsc_0_2_AWLOCK,
      twiddle_h_rsc_0_2_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_2_AWBURST,
      twiddle_h_rsc_0_2_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_2_AWSIZE,
      twiddle_h_rsc_0_2_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_2_AWLEN,
      twiddle_h_rsc_0_2_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_2_AWADDR,
      twiddle_h_rsc_0_2_AWID => twiddle_h_rsc_0_2_AWID,
      twiddle_h_rsc_triosy_0_2_lz => twiddle_h_rsc_triosy_0_2_lz,
      twiddle_h_rsc_0_3_s_tdone => twiddle_h_rsc_0_3_s_tdone,
      twiddle_h_rsc_0_3_tr_write_done => twiddle_h_rsc_0_3_tr_write_done,
      twiddle_h_rsc_0_3_RREADY => twiddle_h_rsc_0_3_RREADY,
      twiddle_h_rsc_0_3_RVALID => twiddle_h_rsc_0_3_RVALID,
      twiddle_h_rsc_0_3_RUSER => twiddle_h_rsc_0_3_RUSER,
      twiddle_h_rsc_0_3_RLAST => twiddle_h_rsc_0_3_RLAST,
      twiddle_h_rsc_0_3_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_3_RRESP,
      twiddle_h_rsc_0_3_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_3_RDATA,
      twiddle_h_rsc_0_3_RID => twiddle_h_rsc_0_3_RID,
      twiddle_h_rsc_0_3_ARREADY => twiddle_h_rsc_0_3_ARREADY,
      twiddle_h_rsc_0_3_ARVALID => twiddle_h_rsc_0_3_ARVALID,
      twiddle_h_rsc_0_3_ARUSER => twiddle_h_rsc_0_3_ARUSER,
      twiddle_h_rsc_0_3_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_3_ARREGION,
      twiddle_h_rsc_0_3_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_3_ARQOS,
      twiddle_h_rsc_0_3_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_3_ARPROT,
      twiddle_h_rsc_0_3_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_3_ARCACHE,
      twiddle_h_rsc_0_3_ARLOCK => twiddle_h_rsc_0_3_ARLOCK,
      twiddle_h_rsc_0_3_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_3_ARBURST,
      twiddle_h_rsc_0_3_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_3_ARSIZE,
      twiddle_h_rsc_0_3_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_3_ARLEN,
      twiddle_h_rsc_0_3_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_3_ARADDR,
      twiddle_h_rsc_0_3_ARID => twiddle_h_rsc_0_3_ARID,
      twiddle_h_rsc_0_3_BREADY => twiddle_h_rsc_0_3_BREADY,
      twiddle_h_rsc_0_3_BVALID => twiddle_h_rsc_0_3_BVALID,
      twiddle_h_rsc_0_3_BUSER => twiddle_h_rsc_0_3_BUSER,
      twiddle_h_rsc_0_3_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_3_BRESP,
      twiddle_h_rsc_0_3_BID => twiddle_h_rsc_0_3_BID,
      twiddle_h_rsc_0_3_WREADY => twiddle_h_rsc_0_3_WREADY,
      twiddle_h_rsc_0_3_WVALID => twiddle_h_rsc_0_3_WVALID,
      twiddle_h_rsc_0_3_WUSER => twiddle_h_rsc_0_3_WUSER,
      twiddle_h_rsc_0_3_WLAST => twiddle_h_rsc_0_3_WLAST,
      twiddle_h_rsc_0_3_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_3_WSTRB,
      twiddle_h_rsc_0_3_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_3_WDATA,
      twiddle_h_rsc_0_3_AWREADY => twiddle_h_rsc_0_3_AWREADY,
      twiddle_h_rsc_0_3_AWVALID => twiddle_h_rsc_0_3_AWVALID,
      twiddle_h_rsc_0_3_AWUSER => twiddle_h_rsc_0_3_AWUSER,
      twiddle_h_rsc_0_3_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_3_AWREGION,
      twiddle_h_rsc_0_3_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_3_AWQOS,
      twiddle_h_rsc_0_3_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_3_AWPROT,
      twiddle_h_rsc_0_3_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_3_AWCACHE,
      twiddle_h_rsc_0_3_AWLOCK => twiddle_h_rsc_0_3_AWLOCK,
      twiddle_h_rsc_0_3_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_3_AWBURST,
      twiddle_h_rsc_0_3_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_3_AWSIZE,
      twiddle_h_rsc_0_3_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_3_AWLEN,
      twiddle_h_rsc_0_3_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_3_AWADDR,
      twiddle_h_rsc_0_3_AWID => twiddle_h_rsc_0_3_AWID,
      twiddle_h_rsc_triosy_0_3_lz => twiddle_h_rsc_triosy_0_3_lz,
      twiddle_h_rsc_0_4_s_tdone => twiddle_h_rsc_0_4_s_tdone,
      twiddle_h_rsc_0_4_tr_write_done => twiddle_h_rsc_0_4_tr_write_done,
      twiddle_h_rsc_0_4_RREADY => twiddle_h_rsc_0_4_RREADY,
      twiddle_h_rsc_0_4_RVALID => twiddle_h_rsc_0_4_RVALID,
      twiddle_h_rsc_0_4_RUSER => twiddle_h_rsc_0_4_RUSER,
      twiddle_h_rsc_0_4_RLAST => twiddle_h_rsc_0_4_RLAST,
      twiddle_h_rsc_0_4_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_4_RRESP,
      twiddle_h_rsc_0_4_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_4_RDATA,
      twiddle_h_rsc_0_4_RID => twiddle_h_rsc_0_4_RID,
      twiddle_h_rsc_0_4_ARREADY => twiddle_h_rsc_0_4_ARREADY,
      twiddle_h_rsc_0_4_ARVALID => twiddle_h_rsc_0_4_ARVALID,
      twiddle_h_rsc_0_4_ARUSER => twiddle_h_rsc_0_4_ARUSER,
      twiddle_h_rsc_0_4_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_4_ARREGION,
      twiddle_h_rsc_0_4_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_4_ARQOS,
      twiddle_h_rsc_0_4_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_4_ARPROT,
      twiddle_h_rsc_0_4_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_4_ARCACHE,
      twiddle_h_rsc_0_4_ARLOCK => twiddle_h_rsc_0_4_ARLOCK,
      twiddle_h_rsc_0_4_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_4_ARBURST,
      twiddle_h_rsc_0_4_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_4_ARSIZE,
      twiddle_h_rsc_0_4_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_4_ARLEN,
      twiddle_h_rsc_0_4_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_4_ARADDR,
      twiddle_h_rsc_0_4_ARID => twiddle_h_rsc_0_4_ARID,
      twiddle_h_rsc_0_4_BREADY => twiddle_h_rsc_0_4_BREADY,
      twiddle_h_rsc_0_4_BVALID => twiddle_h_rsc_0_4_BVALID,
      twiddle_h_rsc_0_4_BUSER => twiddle_h_rsc_0_4_BUSER,
      twiddle_h_rsc_0_4_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_4_BRESP,
      twiddle_h_rsc_0_4_BID => twiddle_h_rsc_0_4_BID,
      twiddle_h_rsc_0_4_WREADY => twiddle_h_rsc_0_4_WREADY,
      twiddle_h_rsc_0_4_WVALID => twiddle_h_rsc_0_4_WVALID,
      twiddle_h_rsc_0_4_WUSER => twiddle_h_rsc_0_4_WUSER,
      twiddle_h_rsc_0_4_WLAST => twiddle_h_rsc_0_4_WLAST,
      twiddle_h_rsc_0_4_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_4_WSTRB,
      twiddle_h_rsc_0_4_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_4_WDATA,
      twiddle_h_rsc_0_4_AWREADY => twiddle_h_rsc_0_4_AWREADY,
      twiddle_h_rsc_0_4_AWVALID => twiddle_h_rsc_0_4_AWVALID,
      twiddle_h_rsc_0_4_AWUSER => twiddle_h_rsc_0_4_AWUSER,
      twiddle_h_rsc_0_4_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_4_AWREGION,
      twiddle_h_rsc_0_4_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_4_AWQOS,
      twiddle_h_rsc_0_4_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_4_AWPROT,
      twiddle_h_rsc_0_4_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_4_AWCACHE,
      twiddle_h_rsc_0_4_AWLOCK => twiddle_h_rsc_0_4_AWLOCK,
      twiddle_h_rsc_0_4_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_4_AWBURST,
      twiddle_h_rsc_0_4_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_4_AWSIZE,
      twiddle_h_rsc_0_4_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_4_AWLEN,
      twiddle_h_rsc_0_4_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_4_AWADDR,
      twiddle_h_rsc_0_4_AWID => twiddle_h_rsc_0_4_AWID,
      twiddle_h_rsc_triosy_0_4_lz => twiddle_h_rsc_triosy_0_4_lz,
      twiddle_h_rsc_0_5_s_tdone => twiddle_h_rsc_0_5_s_tdone,
      twiddle_h_rsc_0_5_tr_write_done => twiddle_h_rsc_0_5_tr_write_done,
      twiddle_h_rsc_0_5_RREADY => twiddle_h_rsc_0_5_RREADY,
      twiddle_h_rsc_0_5_RVALID => twiddle_h_rsc_0_5_RVALID,
      twiddle_h_rsc_0_5_RUSER => twiddle_h_rsc_0_5_RUSER,
      twiddle_h_rsc_0_5_RLAST => twiddle_h_rsc_0_5_RLAST,
      twiddle_h_rsc_0_5_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_5_RRESP,
      twiddle_h_rsc_0_5_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_5_RDATA,
      twiddle_h_rsc_0_5_RID => twiddle_h_rsc_0_5_RID,
      twiddle_h_rsc_0_5_ARREADY => twiddle_h_rsc_0_5_ARREADY,
      twiddle_h_rsc_0_5_ARVALID => twiddle_h_rsc_0_5_ARVALID,
      twiddle_h_rsc_0_5_ARUSER => twiddle_h_rsc_0_5_ARUSER,
      twiddle_h_rsc_0_5_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_5_ARREGION,
      twiddle_h_rsc_0_5_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_5_ARQOS,
      twiddle_h_rsc_0_5_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_5_ARPROT,
      twiddle_h_rsc_0_5_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_5_ARCACHE,
      twiddle_h_rsc_0_5_ARLOCK => twiddle_h_rsc_0_5_ARLOCK,
      twiddle_h_rsc_0_5_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_5_ARBURST,
      twiddle_h_rsc_0_5_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_5_ARSIZE,
      twiddle_h_rsc_0_5_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_5_ARLEN,
      twiddle_h_rsc_0_5_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_5_ARADDR,
      twiddle_h_rsc_0_5_ARID => twiddle_h_rsc_0_5_ARID,
      twiddle_h_rsc_0_5_BREADY => twiddle_h_rsc_0_5_BREADY,
      twiddle_h_rsc_0_5_BVALID => twiddle_h_rsc_0_5_BVALID,
      twiddle_h_rsc_0_5_BUSER => twiddle_h_rsc_0_5_BUSER,
      twiddle_h_rsc_0_5_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_5_BRESP,
      twiddle_h_rsc_0_5_BID => twiddle_h_rsc_0_5_BID,
      twiddle_h_rsc_0_5_WREADY => twiddle_h_rsc_0_5_WREADY,
      twiddle_h_rsc_0_5_WVALID => twiddle_h_rsc_0_5_WVALID,
      twiddle_h_rsc_0_5_WUSER => twiddle_h_rsc_0_5_WUSER,
      twiddle_h_rsc_0_5_WLAST => twiddle_h_rsc_0_5_WLAST,
      twiddle_h_rsc_0_5_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_5_WSTRB,
      twiddle_h_rsc_0_5_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_5_WDATA,
      twiddle_h_rsc_0_5_AWREADY => twiddle_h_rsc_0_5_AWREADY,
      twiddle_h_rsc_0_5_AWVALID => twiddle_h_rsc_0_5_AWVALID,
      twiddle_h_rsc_0_5_AWUSER => twiddle_h_rsc_0_5_AWUSER,
      twiddle_h_rsc_0_5_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_5_AWREGION,
      twiddle_h_rsc_0_5_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_5_AWQOS,
      twiddle_h_rsc_0_5_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_5_AWPROT,
      twiddle_h_rsc_0_5_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_5_AWCACHE,
      twiddle_h_rsc_0_5_AWLOCK => twiddle_h_rsc_0_5_AWLOCK,
      twiddle_h_rsc_0_5_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_5_AWBURST,
      twiddle_h_rsc_0_5_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_5_AWSIZE,
      twiddle_h_rsc_0_5_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_5_AWLEN,
      twiddle_h_rsc_0_5_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_5_AWADDR,
      twiddle_h_rsc_0_5_AWID => twiddle_h_rsc_0_5_AWID,
      twiddle_h_rsc_triosy_0_5_lz => twiddle_h_rsc_triosy_0_5_lz,
      twiddle_h_rsc_0_6_s_tdone => twiddle_h_rsc_0_6_s_tdone,
      twiddle_h_rsc_0_6_tr_write_done => twiddle_h_rsc_0_6_tr_write_done,
      twiddle_h_rsc_0_6_RREADY => twiddle_h_rsc_0_6_RREADY,
      twiddle_h_rsc_0_6_RVALID => twiddle_h_rsc_0_6_RVALID,
      twiddle_h_rsc_0_6_RUSER => twiddle_h_rsc_0_6_RUSER,
      twiddle_h_rsc_0_6_RLAST => twiddle_h_rsc_0_6_RLAST,
      twiddle_h_rsc_0_6_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_6_RRESP,
      twiddle_h_rsc_0_6_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_6_RDATA,
      twiddle_h_rsc_0_6_RID => twiddle_h_rsc_0_6_RID,
      twiddle_h_rsc_0_6_ARREADY => twiddle_h_rsc_0_6_ARREADY,
      twiddle_h_rsc_0_6_ARVALID => twiddle_h_rsc_0_6_ARVALID,
      twiddle_h_rsc_0_6_ARUSER => twiddle_h_rsc_0_6_ARUSER,
      twiddle_h_rsc_0_6_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_6_ARREGION,
      twiddle_h_rsc_0_6_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_6_ARQOS,
      twiddle_h_rsc_0_6_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_6_ARPROT,
      twiddle_h_rsc_0_6_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_6_ARCACHE,
      twiddle_h_rsc_0_6_ARLOCK => twiddle_h_rsc_0_6_ARLOCK,
      twiddle_h_rsc_0_6_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_6_ARBURST,
      twiddle_h_rsc_0_6_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_6_ARSIZE,
      twiddle_h_rsc_0_6_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_6_ARLEN,
      twiddle_h_rsc_0_6_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_6_ARADDR,
      twiddle_h_rsc_0_6_ARID => twiddle_h_rsc_0_6_ARID,
      twiddle_h_rsc_0_6_BREADY => twiddle_h_rsc_0_6_BREADY,
      twiddle_h_rsc_0_6_BVALID => twiddle_h_rsc_0_6_BVALID,
      twiddle_h_rsc_0_6_BUSER => twiddle_h_rsc_0_6_BUSER,
      twiddle_h_rsc_0_6_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_6_BRESP,
      twiddle_h_rsc_0_6_BID => twiddle_h_rsc_0_6_BID,
      twiddle_h_rsc_0_6_WREADY => twiddle_h_rsc_0_6_WREADY,
      twiddle_h_rsc_0_6_WVALID => twiddle_h_rsc_0_6_WVALID,
      twiddle_h_rsc_0_6_WUSER => twiddle_h_rsc_0_6_WUSER,
      twiddle_h_rsc_0_6_WLAST => twiddle_h_rsc_0_6_WLAST,
      twiddle_h_rsc_0_6_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_6_WSTRB,
      twiddle_h_rsc_0_6_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_6_WDATA,
      twiddle_h_rsc_0_6_AWREADY => twiddle_h_rsc_0_6_AWREADY,
      twiddle_h_rsc_0_6_AWVALID => twiddle_h_rsc_0_6_AWVALID,
      twiddle_h_rsc_0_6_AWUSER => twiddle_h_rsc_0_6_AWUSER,
      twiddle_h_rsc_0_6_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_6_AWREGION,
      twiddle_h_rsc_0_6_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_6_AWQOS,
      twiddle_h_rsc_0_6_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_6_AWPROT,
      twiddle_h_rsc_0_6_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_6_AWCACHE,
      twiddle_h_rsc_0_6_AWLOCK => twiddle_h_rsc_0_6_AWLOCK,
      twiddle_h_rsc_0_6_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_6_AWBURST,
      twiddle_h_rsc_0_6_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_6_AWSIZE,
      twiddle_h_rsc_0_6_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_6_AWLEN,
      twiddle_h_rsc_0_6_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_6_AWADDR,
      twiddle_h_rsc_0_6_AWID => twiddle_h_rsc_0_6_AWID,
      twiddle_h_rsc_triosy_0_6_lz => twiddle_h_rsc_triosy_0_6_lz,
      twiddle_h_rsc_0_7_s_tdone => twiddle_h_rsc_0_7_s_tdone,
      twiddle_h_rsc_0_7_tr_write_done => twiddle_h_rsc_0_7_tr_write_done,
      twiddle_h_rsc_0_7_RREADY => twiddle_h_rsc_0_7_RREADY,
      twiddle_h_rsc_0_7_RVALID => twiddle_h_rsc_0_7_RVALID,
      twiddle_h_rsc_0_7_RUSER => twiddle_h_rsc_0_7_RUSER,
      twiddle_h_rsc_0_7_RLAST => twiddle_h_rsc_0_7_RLAST,
      twiddle_h_rsc_0_7_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_7_RRESP,
      twiddle_h_rsc_0_7_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_7_RDATA,
      twiddle_h_rsc_0_7_RID => twiddle_h_rsc_0_7_RID,
      twiddle_h_rsc_0_7_ARREADY => twiddle_h_rsc_0_7_ARREADY,
      twiddle_h_rsc_0_7_ARVALID => twiddle_h_rsc_0_7_ARVALID,
      twiddle_h_rsc_0_7_ARUSER => twiddle_h_rsc_0_7_ARUSER,
      twiddle_h_rsc_0_7_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_7_ARREGION,
      twiddle_h_rsc_0_7_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_7_ARQOS,
      twiddle_h_rsc_0_7_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_7_ARPROT,
      twiddle_h_rsc_0_7_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_7_ARCACHE,
      twiddle_h_rsc_0_7_ARLOCK => twiddle_h_rsc_0_7_ARLOCK,
      twiddle_h_rsc_0_7_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_7_ARBURST,
      twiddle_h_rsc_0_7_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_7_ARSIZE,
      twiddle_h_rsc_0_7_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_7_ARLEN,
      twiddle_h_rsc_0_7_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_7_ARADDR,
      twiddle_h_rsc_0_7_ARID => twiddle_h_rsc_0_7_ARID,
      twiddle_h_rsc_0_7_BREADY => twiddle_h_rsc_0_7_BREADY,
      twiddle_h_rsc_0_7_BVALID => twiddle_h_rsc_0_7_BVALID,
      twiddle_h_rsc_0_7_BUSER => twiddle_h_rsc_0_7_BUSER,
      twiddle_h_rsc_0_7_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_7_BRESP,
      twiddle_h_rsc_0_7_BID => twiddle_h_rsc_0_7_BID,
      twiddle_h_rsc_0_7_WREADY => twiddle_h_rsc_0_7_WREADY,
      twiddle_h_rsc_0_7_WVALID => twiddle_h_rsc_0_7_WVALID,
      twiddle_h_rsc_0_7_WUSER => twiddle_h_rsc_0_7_WUSER,
      twiddle_h_rsc_0_7_WLAST => twiddle_h_rsc_0_7_WLAST,
      twiddle_h_rsc_0_7_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_7_WSTRB,
      twiddle_h_rsc_0_7_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_7_WDATA,
      twiddle_h_rsc_0_7_AWREADY => twiddle_h_rsc_0_7_AWREADY,
      twiddle_h_rsc_0_7_AWVALID => twiddle_h_rsc_0_7_AWVALID,
      twiddle_h_rsc_0_7_AWUSER => twiddle_h_rsc_0_7_AWUSER,
      twiddle_h_rsc_0_7_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_7_AWREGION,
      twiddle_h_rsc_0_7_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_7_AWQOS,
      twiddle_h_rsc_0_7_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_7_AWPROT,
      twiddle_h_rsc_0_7_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_7_AWCACHE,
      twiddle_h_rsc_0_7_AWLOCK => twiddle_h_rsc_0_7_AWLOCK,
      twiddle_h_rsc_0_7_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_7_AWBURST,
      twiddle_h_rsc_0_7_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_7_AWSIZE,
      twiddle_h_rsc_0_7_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_7_AWLEN,
      twiddle_h_rsc_0_7_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_7_AWADDR,
      twiddle_h_rsc_0_7_AWID => twiddle_h_rsc_0_7_AWID,
      twiddle_h_rsc_triosy_0_7_lz => twiddle_h_rsc_triosy_0_7_lz,
      twiddle_h_rsc_0_8_s_tdone => twiddle_h_rsc_0_8_s_tdone,
      twiddle_h_rsc_0_8_tr_write_done => twiddle_h_rsc_0_8_tr_write_done,
      twiddle_h_rsc_0_8_RREADY => twiddle_h_rsc_0_8_RREADY,
      twiddle_h_rsc_0_8_RVALID => twiddle_h_rsc_0_8_RVALID,
      twiddle_h_rsc_0_8_RUSER => twiddle_h_rsc_0_8_RUSER,
      twiddle_h_rsc_0_8_RLAST => twiddle_h_rsc_0_8_RLAST,
      twiddle_h_rsc_0_8_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_8_RRESP,
      twiddle_h_rsc_0_8_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_8_RDATA,
      twiddle_h_rsc_0_8_RID => twiddle_h_rsc_0_8_RID,
      twiddle_h_rsc_0_8_ARREADY => twiddle_h_rsc_0_8_ARREADY,
      twiddle_h_rsc_0_8_ARVALID => twiddle_h_rsc_0_8_ARVALID,
      twiddle_h_rsc_0_8_ARUSER => twiddle_h_rsc_0_8_ARUSER,
      twiddle_h_rsc_0_8_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_8_ARREGION,
      twiddle_h_rsc_0_8_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_8_ARQOS,
      twiddle_h_rsc_0_8_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_8_ARPROT,
      twiddle_h_rsc_0_8_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_8_ARCACHE,
      twiddle_h_rsc_0_8_ARLOCK => twiddle_h_rsc_0_8_ARLOCK,
      twiddle_h_rsc_0_8_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_8_ARBURST,
      twiddle_h_rsc_0_8_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_8_ARSIZE,
      twiddle_h_rsc_0_8_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_8_ARLEN,
      twiddle_h_rsc_0_8_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_8_ARADDR,
      twiddle_h_rsc_0_8_ARID => twiddle_h_rsc_0_8_ARID,
      twiddle_h_rsc_0_8_BREADY => twiddle_h_rsc_0_8_BREADY,
      twiddle_h_rsc_0_8_BVALID => twiddle_h_rsc_0_8_BVALID,
      twiddle_h_rsc_0_8_BUSER => twiddle_h_rsc_0_8_BUSER,
      twiddle_h_rsc_0_8_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_8_BRESP,
      twiddle_h_rsc_0_8_BID => twiddle_h_rsc_0_8_BID,
      twiddle_h_rsc_0_8_WREADY => twiddle_h_rsc_0_8_WREADY,
      twiddle_h_rsc_0_8_WVALID => twiddle_h_rsc_0_8_WVALID,
      twiddle_h_rsc_0_8_WUSER => twiddle_h_rsc_0_8_WUSER,
      twiddle_h_rsc_0_8_WLAST => twiddle_h_rsc_0_8_WLAST,
      twiddle_h_rsc_0_8_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_8_WSTRB,
      twiddle_h_rsc_0_8_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_8_WDATA,
      twiddle_h_rsc_0_8_AWREADY => twiddle_h_rsc_0_8_AWREADY,
      twiddle_h_rsc_0_8_AWVALID => twiddle_h_rsc_0_8_AWVALID,
      twiddle_h_rsc_0_8_AWUSER => twiddle_h_rsc_0_8_AWUSER,
      twiddle_h_rsc_0_8_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_8_AWREGION,
      twiddle_h_rsc_0_8_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_8_AWQOS,
      twiddle_h_rsc_0_8_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_8_AWPROT,
      twiddle_h_rsc_0_8_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_8_AWCACHE,
      twiddle_h_rsc_0_8_AWLOCK => twiddle_h_rsc_0_8_AWLOCK,
      twiddle_h_rsc_0_8_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_8_AWBURST,
      twiddle_h_rsc_0_8_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_8_AWSIZE,
      twiddle_h_rsc_0_8_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_8_AWLEN,
      twiddle_h_rsc_0_8_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_8_AWADDR,
      twiddle_h_rsc_0_8_AWID => twiddle_h_rsc_0_8_AWID,
      twiddle_h_rsc_triosy_0_8_lz => twiddle_h_rsc_triosy_0_8_lz,
      twiddle_h_rsc_0_9_s_tdone => twiddle_h_rsc_0_9_s_tdone,
      twiddle_h_rsc_0_9_tr_write_done => twiddle_h_rsc_0_9_tr_write_done,
      twiddle_h_rsc_0_9_RREADY => twiddle_h_rsc_0_9_RREADY,
      twiddle_h_rsc_0_9_RVALID => twiddle_h_rsc_0_9_RVALID,
      twiddle_h_rsc_0_9_RUSER => twiddle_h_rsc_0_9_RUSER,
      twiddle_h_rsc_0_9_RLAST => twiddle_h_rsc_0_9_RLAST,
      twiddle_h_rsc_0_9_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_9_RRESP,
      twiddle_h_rsc_0_9_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_9_RDATA,
      twiddle_h_rsc_0_9_RID => twiddle_h_rsc_0_9_RID,
      twiddle_h_rsc_0_9_ARREADY => twiddle_h_rsc_0_9_ARREADY,
      twiddle_h_rsc_0_9_ARVALID => twiddle_h_rsc_0_9_ARVALID,
      twiddle_h_rsc_0_9_ARUSER => twiddle_h_rsc_0_9_ARUSER,
      twiddle_h_rsc_0_9_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_9_ARREGION,
      twiddle_h_rsc_0_9_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_9_ARQOS,
      twiddle_h_rsc_0_9_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_9_ARPROT,
      twiddle_h_rsc_0_9_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_9_ARCACHE,
      twiddle_h_rsc_0_9_ARLOCK => twiddle_h_rsc_0_9_ARLOCK,
      twiddle_h_rsc_0_9_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_9_ARBURST,
      twiddle_h_rsc_0_9_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_9_ARSIZE,
      twiddle_h_rsc_0_9_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_9_ARLEN,
      twiddle_h_rsc_0_9_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_9_ARADDR,
      twiddle_h_rsc_0_9_ARID => twiddle_h_rsc_0_9_ARID,
      twiddle_h_rsc_0_9_BREADY => twiddle_h_rsc_0_9_BREADY,
      twiddle_h_rsc_0_9_BVALID => twiddle_h_rsc_0_9_BVALID,
      twiddle_h_rsc_0_9_BUSER => twiddle_h_rsc_0_9_BUSER,
      twiddle_h_rsc_0_9_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_9_BRESP,
      twiddle_h_rsc_0_9_BID => twiddle_h_rsc_0_9_BID,
      twiddle_h_rsc_0_9_WREADY => twiddle_h_rsc_0_9_WREADY,
      twiddle_h_rsc_0_9_WVALID => twiddle_h_rsc_0_9_WVALID,
      twiddle_h_rsc_0_9_WUSER => twiddle_h_rsc_0_9_WUSER,
      twiddle_h_rsc_0_9_WLAST => twiddle_h_rsc_0_9_WLAST,
      twiddle_h_rsc_0_9_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_9_WSTRB,
      twiddle_h_rsc_0_9_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_9_WDATA,
      twiddle_h_rsc_0_9_AWREADY => twiddle_h_rsc_0_9_AWREADY,
      twiddle_h_rsc_0_9_AWVALID => twiddle_h_rsc_0_9_AWVALID,
      twiddle_h_rsc_0_9_AWUSER => twiddle_h_rsc_0_9_AWUSER,
      twiddle_h_rsc_0_9_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_9_AWREGION,
      twiddle_h_rsc_0_9_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_9_AWQOS,
      twiddle_h_rsc_0_9_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_9_AWPROT,
      twiddle_h_rsc_0_9_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_9_AWCACHE,
      twiddle_h_rsc_0_9_AWLOCK => twiddle_h_rsc_0_9_AWLOCK,
      twiddle_h_rsc_0_9_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_9_AWBURST,
      twiddle_h_rsc_0_9_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_9_AWSIZE,
      twiddle_h_rsc_0_9_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_9_AWLEN,
      twiddle_h_rsc_0_9_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_9_AWADDR,
      twiddle_h_rsc_0_9_AWID => twiddle_h_rsc_0_9_AWID,
      twiddle_h_rsc_triosy_0_9_lz => twiddle_h_rsc_triosy_0_9_lz,
      twiddle_h_rsc_0_10_s_tdone => twiddle_h_rsc_0_10_s_tdone,
      twiddle_h_rsc_0_10_tr_write_done => twiddle_h_rsc_0_10_tr_write_done,
      twiddle_h_rsc_0_10_RREADY => twiddle_h_rsc_0_10_RREADY,
      twiddle_h_rsc_0_10_RVALID => twiddle_h_rsc_0_10_RVALID,
      twiddle_h_rsc_0_10_RUSER => twiddle_h_rsc_0_10_RUSER,
      twiddle_h_rsc_0_10_RLAST => twiddle_h_rsc_0_10_RLAST,
      twiddle_h_rsc_0_10_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_10_RRESP,
      twiddle_h_rsc_0_10_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_10_RDATA,
      twiddle_h_rsc_0_10_RID => twiddle_h_rsc_0_10_RID,
      twiddle_h_rsc_0_10_ARREADY => twiddle_h_rsc_0_10_ARREADY,
      twiddle_h_rsc_0_10_ARVALID => twiddle_h_rsc_0_10_ARVALID,
      twiddle_h_rsc_0_10_ARUSER => twiddle_h_rsc_0_10_ARUSER,
      twiddle_h_rsc_0_10_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_10_ARREGION,
      twiddle_h_rsc_0_10_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_10_ARQOS,
      twiddle_h_rsc_0_10_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_10_ARPROT,
      twiddle_h_rsc_0_10_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_10_ARCACHE,
      twiddle_h_rsc_0_10_ARLOCK => twiddle_h_rsc_0_10_ARLOCK,
      twiddle_h_rsc_0_10_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_10_ARBURST,
      twiddle_h_rsc_0_10_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_10_ARSIZE,
      twiddle_h_rsc_0_10_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_10_ARLEN,
      twiddle_h_rsc_0_10_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_10_ARADDR,
      twiddle_h_rsc_0_10_ARID => twiddle_h_rsc_0_10_ARID,
      twiddle_h_rsc_0_10_BREADY => twiddle_h_rsc_0_10_BREADY,
      twiddle_h_rsc_0_10_BVALID => twiddle_h_rsc_0_10_BVALID,
      twiddle_h_rsc_0_10_BUSER => twiddle_h_rsc_0_10_BUSER,
      twiddle_h_rsc_0_10_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_10_BRESP,
      twiddle_h_rsc_0_10_BID => twiddle_h_rsc_0_10_BID,
      twiddle_h_rsc_0_10_WREADY => twiddle_h_rsc_0_10_WREADY,
      twiddle_h_rsc_0_10_WVALID => twiddle_h_rsc_0_10_WVALID,
      twiddle_h_rsc_0_10_WUSER => twiddle_h_rsc_0_10_WUSER,
      twiddle_h_rsc_0_10_WLAST => twiddle_h_rsc_0_10_WLAST,
      twiddle_h_rsc_0_10_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_10_WSTRB,
      twiddle_h_rsc_0_10_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_10_WDATA,
      twiddle_h_rsc_0_10_AWREADY => twiddle_h_rsc_0_10_AWREADY,
      twiddle_h_rsc_0_10_AWVALID => twiddle_h_rsc_0_10_AWVALID,
      twiddle_h_rsc_0_10_AWUSER => twiddle_h_rsc_0_10_AWUSER,
      twiddle_h_rsc_0_10_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_10_AWREGION,
      twiddle_h_rsc_0_10_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_10_AWQOS,
      twiddle_h_rsc_0_10_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_10_AWPROT,
      twiddle_h_rsc_0_10_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_10_AWCACHE,
      twiddle_h_rsc_0_10_AWLOCK => twiddle_h_rsc_0_10_AWLOCK,
      twiddle_h_rsc_0_10_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_10_AWBURST,
      twiddle_h_rsc_0_10_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_10_AWSIZE,
      twiddle_h_rsc_0_10_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_10_AWLEN,
      twiddle_h_rsc_0_10_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_10_AWADDR,
      twiddle_h_rsc_0_10_AWID => twiddle_h_rsc_0_10_AWID,
      twiddle_h_rsc_triosy_0_10_lz => twiddle_h_rsc_triosy_0_10_lz,
      twiddle_h_rsc_0_11_s_tdone => twiddle_h_rsc_0_11_s_tdone,
      twiddle_h_rsc_0_11_tr_write_done => twiddle_h_rsc_0_11_tr_write_done,
      twiddle_h_rsc_0_11_RREADY => twiddle_h_rsc_0_11_RREADY,
      twiddle_h_rsc_0_11_RVALID => twiddle_h_rsc_0_11_RVALID,
      twiddle_h_rsc_0_11_RUSER => twiddle_h_rsc_0_11_RUSER,
      twiddle_h_rsc_0_11_RLAST => twiddle_h_rsc_0_11_RLAST,
      twiddle_h_rsc_0_11_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_11_RRESP,
      twiddle_h_rsc_0_11_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_11_RDATA,
      twiddle_h_rsc_0_11_RID => twiddle_h_rsc_0_11_RID,
      twiddle_h_rsc_0_11_ARREADY => twiddle_h_rsc_0_11_ARREADY,
      twiddle_h_rsc_0_11_ARVALID => twiddle_h_rsc_0_11_ARVALID,
      twiddle_h_rsc_0_11_ARUSER => twiddle_h_rsc_0_11_ARUSER,
      twiddle_h_rsc_0_11_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_11_ARREGION,
      twiddle_h_rsc_0_11_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_11_ARQOS,
      twiddle_h_rsc_0_11_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_11_ARPROT,
      twiddle_h_rsc_0_11_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_11_ARCACHE,
      twiddle_h_rsc_0_11_ARLOCK => twiddle_h_rsc_0_11_ARLOCK,
      twiddle_h_rsc_0_11_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_11_ARBURST,
      twiddle_h_rsc_0_11_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_11_ARSIZE,
      twiddle_h_rsc_0_11_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_11_ARLEN,
      twiddle_h_rsc_0_11_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_11_ARADDR,
      twiddle_h_rsc_0_11_ARID => twiddle_h_rsc_0_11_ARID,
      twiddle_h_rsc_0_11_BREADY => twiddle_h_rsc_0_11_BREADY,
      twiddle_h_rsc_0_11_BVALID => twiddle_h_rsc_0_11_BVALID,
      twiddle_h_rsc_0_11_BUSER => twiddle_h_rsc_0_11_BUSER,
      twiddle_h_rsc_0_11_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_11_BRESP,
      twiddle_h_rsc_0_11_BID => twiddle_h_rsc_0_11_BID,
      twiddle_h_rsc_0_11_WREADY => twiddle_h_rsc_0_11_WREADY,
      twiddle_h_rsc_0_11_WVALID => twiddle_h_rsc_0_11_WVALID,
      twiddle_h_rsc_0_11_WUSER => twiddle_h_rsc_0_11_WUSER,
      twiddle_h_rsc_0_11_WLAST => twiddle_h_rsc_0_11_WLAST,
      twiddle_h_rsc_0_11_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_11_WSTRB,
      twiddle_h_rsc_0_11_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_11_WDATA,
      twiddle_h_rsc_0_11_AWREADY => twiddle_h_rsc_0_11_AWREADY,
      twiddle_h_rsc_0_11_AWVALID => twiddle_h_rsc_0_11_AWVALID,
      twiddle_h_rsc_0_11_AWUSER => twiddle_h_rsc_0_11_AWUSER,
      twiddle_h_rsc_0_11_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_11_AWREGION,
      twiddle_h_rsc_0_11_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_11_AWQOS,
      twiddle_h_rsc_0_11_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_11_AWPROT,
      twiddle_h_rsc_0_11_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_11_AWCACHE,
      twiddle_h_rsc_0_11_AWLOCK => twiddle_h_rsc_0_11_AWLOCK,
      twiddle_h_rsc_0_11_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_11_AWBURST,
      twiddle_h_rsc_0_11_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_11_AWSIZE,
      twiddle_h_rsc_0_11_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_11_AWLEN,
      twiddle_h_rsc_0_11_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_11_AWADDR,
      twiddle_h_rsc_0_11_AWID => twiddle_h_rsc_0_11_AWID,
      twiddle_h_rsc_triosy_0_11_lz => twiddle_h_rsc_triosy_0_11_lz,
      twiddle_h_rsc_0_12_s_tdone => twiddle_h_rsc_0_12_s_tdone,
      twiddle_h_rsc_0_12_tr_write_done => twiddle_h_rsc_0_12_tr_write_done,
      twiddle_h_rsc_0_12_RREADY => twiddle_h_rsc_0_12_RREADY,
      twiddle_h_rsc_0_12_RVALID => twiddle_h_rsc_0_12_RVALID,
      twiddle_h_rsc_0_12_RUSER => twiddle_h_rsc_0_12_RUSER,
      twiddle_h_rsc_0_12_RLAST => twiddle_h_rsc_0_12_RLAST,
      twiddle_h_rsc_0_12_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_12_RRESP,
      twiddle_h_rsc_0_12_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_12_RDATA,
      twiddle_h_rsc_0_12_RID => twiddle_h_rsc_0_12_RID,
      twiddle_h_rsc_0_12_ARREADY => twiddle_h_rsc_0_12_ARREADY,
      twiddle_h_rsc_0_12_ARVALID => twiddle_h_rsc_0_12_ARVALID,
      twiddle_h_rsc_0_12_ARUSER => twiddle_h_rsc_0_12_ARUSER,
      twiddle_h_rsc_0_12_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_12_ARREGION,
      twiddle_h_rsc_0_12_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_12_ARQOS,
      twiddle_h_rsc_0_12_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_12_ARPROT,
      twiddle_h_rsc_0_12_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_12_ARCACHE,
      twiddle_h_rsc_0_12_ARLOCK => twiddle_h_rsc_0_12_ARLOCK,
      twiddle_h_rsc_0_12_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_12_ARBURST,
      twiddle_h_rsc_0_12_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_12_ARSIZE,
      twiddle_h_rsc_0_12_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_12_ARLEN,
      twiddle_h_rsc_0_12_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_12_ARADDR,
      twiddle_h_rsc_0_12_ARID => twiddle_h_rsc_0_12_ARID,
      twiddle_h_rsc_0_12_BREADY => twiddle_h_rsc_0_12_BREADY,
      twiddle_h_rsc_0_12_BVALID => twiddle_h_rsc_0_12_BVALID,
      twiddle_h_rsc_0_12_BUSER => twiddle_h_rsc_0_12_BUSER,
      twiddle_h_rsc_0_12_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_12_BRESP,
      twiddle_h_rsc_0_12_BID => twiddle_h_rsc_0_12_BID,
      twiddle_h_rsc_0_12_WREADY => twiddle_h_rsc_0_12_WREADY,
      twiddle_h_rsc_0_12_WVALID => twiddle_h_rsc_0_12_WVALID,
      twiddle_h_rsc_0_12_WUSER => twiddle_h_rsc_0_12_WUSER,
      twiddle_h_rsc_0_12_WLAST => twiddle_h_rsc_0_12_WLAST,
      twiddle_h_rsc_0_12_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_12_WSTRB,
      twiddle_h_rsc_0_12_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_12_WDATA,
      twiddle_h_rsc_0_12_AWREADY => twiddle_h_rsc_0_12_AWREADY,
      twiddle_h_rsc_0_12_AWVALID => twiddle_h_rsc_0_12_AWVALID,
      twiddle_h_rsc_0_12_AWUSER => twiddle_h_rsc_0_12_AWUSER,
      twiddle_h_rsc_0_12_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_12_AWREGION,
      twiddle_h_rsc_0_12_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_12_AWQOS,
      twiddle_h_rsc_0_12_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_12_AWPROT,
      twiddle_h_rsc_0_12_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_12_AWCACHE,
      twiddle_h_rsc_0_12_AWLOCK => twiddle_h_rsc_0_12_AWLOCK,
      twiddle_h_rsc_0_12_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_12_AWBURST,
      twiddle_h_rsc_0_12_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_12_AWSIZE,
      twiddle_h_rsc_0_12_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_12_AWLEN,
      twiddle_h_rsc_0_12_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_12_AWADDR,
      twiddle_h_rsc_0_12_AWID => twiddle_h_rsc_0_12_AWID,
      twiddle_h_rsc_triosy_0_12_lz => twiddle_h_rsc_triosy_0_12_lz,
      twiddle_h_rsc_0_13_s_tdone => twiddle_h_rsc_0_13_s_tdone,
      twiddle_h_rsc_0_13_tr_write_done => twiddle_h_rsc_0_13_tr_write_done,
      twiddle_h_rsc_0_13_RREADY => twiddle_h_rsc_0_13_RREADY,
      twiddle_h_rsc_0_13_RVALID => twiddle_h_rsc_0_13_RVALID,
      twiddle_h_rsc_0_13_RUSER => twiddle_h_rsc_0_13_RUSER,
      twiddle_h_rsc_0_13_RLAST => twiddle_h_rsc_0_13_RLAST,
      twiddle_h_rsc_0_13_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_13_RRESP,
      twiddle_h_rsc_0_13_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_13_RDATA,
      twiddle_h_rsc_0_13_RID => twiddle_h_rsc_0_13_RID,
      twiddle_h_rsc_0_13_ARREADY => twiddle_h_rsc_0_13_ARREADY,
      twiddle_h_rsc_0_13_ARVALID => twiddle_h_rsc_0_13_ARVALID,
      twiddle_h_rsc_0_13_ARUSER => twiddle_h_rsc_0_13_ARUSER,
      twiddle_h_rsc_0_13_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_13_ARREGION,
      twiddle_h_rsc_0_13_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_13_ARQOS,
      twiddle_h_rsc_0_13_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_13_ARPROT,
      twiddle_h_rsc_0_13_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_13_ARCACHE,
      twiddle_h_rsc_0_13_ARLOCK => twiddle_h_rsc_0_13_ARLOCK,
      twiddle_h_rsc_0_13_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_13_ARBURST,
      twiddle_h_rsc_0_13_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_13_ARSIZE,
      twiddle_h_rsc_0_13_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_13_ARLEN,
      twiddle_h_rsc_0_13_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_13_ARADDR,
      twiddle_h_rsc_0_13_ARID => twiddle_h_rsc_0_13_ARID,
      twiddle_h_rsc_0_13_BREADY => twiddle_h_rsc_0_13_BREADY,
      twiddle_h_rsc_0_13_BVALID => twiddle_h_rsc_0_13_BVALID,
      twiddle_h_rsc_0_13_BUSER => twiddle_h_rsc_0_13_BUSER,
      twiddle_h_rsc_0_13_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_13_BRESP,
      twiddle_h_rsc_0_13_BID => twiddle_h_rsc_0_13_BID,
      twiddle_h_rsc_0_13_WREADY => twiddle_h_rsc_0_13_WREADY,
      twiddle_h_rsc_0_13_WVALID => twiddle_h_rsc_0_13_WVALID,
      twiddle_h_rsc_0_13_WUSER => twiddle_h_rsc_0_13_WUSER,
      twiddle_h_rsc_0_13_WLAST => twiddle_h_rsc_0_13_WLAST,
      twiddle_h_rsc_0_13_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_13_WSTRB,
      twiddle_h_rsc_0_13_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_13_WDATA,
      twiddle_h_rsc_0_13_AWREADY => twiddle_h_rsc_0_13_AWREADY,
      twiddle_h_rsc_0_13_AWVALID => twiddle_h_rsc_0_13_AWVALID,
      twiddle_h_rsc_0_13_AWUSER => twiddle_h_rsc_0_13_AWUSER,
      twiddle_h_rsc_0_13_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_13_AWREGION,
      twiddle_h_rsc_0_13_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_13_AWQOS,
      twiddle_h_rsc_0_13_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_13_AWPROT,
      twiddle_h_rsc_0_13_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_13_AWCACHE,
      twiddle_h_rsc_0_13_AWLOCK => twiddle_h_rsc_0_13_AWLOCK,
      twiddle_h_rsc_0_13_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_13_AWBURST,
      twiddle_h_rsc_0_13_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_13_AWSIZE,
      twiddle_h_rsc_0_13_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_13_AWLEN,
      twiddle_h_rsc_0_13_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_13_AWADDR,
      twiddle_h_rsc_0_13_AWID => twiddle_h_rsc_0_13_AWID,
      twiddle_h_rsc_triosy_0_13_lz => twiddle_h_rsc_triosy_0_13_lz,
      twiddle_h_rsc_0_14_s_tdone => twiddle_h_rsc_0_14_s_tdone,
      twiddle_h_rsc_0_14_tr_write_done => twiddle_h_rsc_0_14_tr_write_done,
      twiddle_h_rsc_0_14_RREADY => twiddle_h_rsc_0_14_RREADY,
      twiddle_h_rsc_0_14_RVALID => twiddle_h_rsc_0_14_RVALID,
      twiddle_h_rsc_0_14_RUSER => twiddle_h_rsc_0_14_RUSER,
      twiddle_h_rsc_0_14_RLAST => twiddle_h_rsc_0_14_RLAST,
      twiddle_h_rsc_0_14_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_14_RRESP,
      twiddle_h_rsc_0_14_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_14_RDATA,
      twiddle_h_rsc_0_14_RID => twiddle_h_rsc_0_14_RID,
      twiddle_h_rsc_0_14_ARREADY => twiddle_h_rsc_0_14_ARREADY,
      twiddle_h_rsc_0_14_ARVALID => twiddle_h_rsc_0_14_ARVALID,
      twiddle_h_rsc_0_14_ARUSER => twiddle_h_rsc_0_14_ARUSER,
      twiddle_h_rsc_0_14_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_14_ARREGION,
      twiddle_h_rsc_0_14_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_14_ARQOS,
      twiddle_h_rsc_0_14_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_14_ARPROT,
      twiddle_h_rsc_0_14_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_14_ARCACHE,
      twiddle_h_rsc_0_14_ARLOCK => twiddle_h_rsc_0_14_ARLOCK,
      twiddle_h_rsc_0_14_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_14_ARBURST,
      twiddle_h_rsc_0_14_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_14_ARSIZE,
      twiddle_h_rsc_0_14_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_14_ARLEN,
      twiddle_h_rsc_0_14_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_14_ARADDR,
      twiddle_h_rsc_0_14_ARID => twiddle_h_rsc_0_14_ARID,
      twiddle_h_rsc_0_14_BREADY => twiddle_h_rsc_0_14_BREADY,
      twiddle_h_rsc_0_14_BVALID => twiddle_h_rsc_0_14_BVALID,
      twiddle_h_rsc_0_14_BUSER => twiddle_h_rsc_0_14_BUSER,
      twiddle_h_rsc_0_14_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_14_BRESP,
      twiddle_h_rsc_0_14_BID => twiddle_h_rsc_0_14_BID,
      twiddle_h_rsc_0_14_WREADY => twiddle_h_rsc_0_14_WREADY,
      twiddle_h_rsc_0_14_WVALID => twiddle_h_rsc_0_14_WVALID,
      twiddle_h_rsc_0_14_WUSER => twiddle_h_rsc_0_14_WUSER,
      twiddle_h_rsc_0_14_WLAST => twiddle_h_rsc_0_14_WLAST,
      twiddle_h_rsc_0_14_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_14_WSTRB,
      twiddle_h_rsc_0_14_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_14_WDATA,
      twiddle_h_rsc_0_14_AWREADY => twiddle_h_rsc_0_14_AWREADY,
      twiddle_h_rsc_0_14_AWVALID => twiddle_h_rsc_0_14_AWVALID,
      twiddle_h_rsc_0_14_AWUSER => twiddle_h_rsc_0_14_AWUSER,
      twiddle_h_rsc_0_14_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_14_AWREGION,
      twiddle_h_rsc_0_14_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_14_AWQOS,
      twiddle_h_rsc_0_14_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_14_AWPROT,
      twiddle_h_rsc_0_14_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_14_AWCACHE,
      twiddle_h_rsc_0_14_AWLOCK => twiddle_h_rsc_0_14_AWLOCK,
      twiddle_h_rsc_0_14_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_14_AWBURST,
      twiddle_h_rsc_0_14_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_14_AWSIZE,
      twiddle_h_rsc_0_14_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_14_AWLEN,
      twiddle_h_rsc_0_14_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_14_AWADDR,
      twiddle_h_rsc_0_14_AWID => twiddle_h_rsc_0_14_AWID,
      twiddle_h_rsc_triosy_0_14_lz => twiddle_h_rsc_triosy_0_14_lz,
      twiddle_h_rsc_0_15_s_tdone => twiddle_h_rsc_0_15_s_tdone,
      twiddle_h_rsc_0_15_tr_write_done => twiddle_h_rsc_0_15_tr_write_done,
      twiddle_h_rsc_0_15_RREADY => twiddle_h_rsc_0_15_RREADY,
      twiddle_h_rsc_0_15_RVALID => twiddle_h_rsc_0_15_RVALID,
      twiddle_h_rsc_0_15_RUSER => twiddle_h_rsc_0_15_RUSER,
      twiddle_h_rsc_0_15_RLAST => twiddle_h_rsc_0_15_RLAST,
      twiddle_h_rsc_0_15_RRESP => peaseNTT_core_inst_twiddle_h_rsc_0_15_RRESP,
      twiddle_h_rsc_0_15_RDATA => peaseNTT_core_inst_twiddle_h_rsc_0_15_RDATA,
      twiddle_h_rsc_0_15_RID => twiddle_h_rsc_0_15_RID,
      twiddle_h_rsc_0_15_ARREADY => twiddle_h_rsc_0_15_ARREADY,
      twiddle_h_rsc_0_15_ARVALID => twiddle_h_rsc_0_15_ARVALID,
      twiddle_h_rsc_0_15_ARUSER => twiddle_h_rsc_0_15_ARUSER,
      twiddle_h_rsc_0_15_ARREGION => peaseNTT_core_inst_twiddle_h_rsc_0_15_ARREGION,
      twiddle_h_rsc_0_15_ARQOS => peaseNTT_core_inst_twiddle_h_rsc_0_15_ARQOS,
      twiddle_h_rsc_0_15_ARPROT => peaseNTT_core_inst_twiddle_h_rsc_0_15_ARPROT,
      twiddle_h_rsc_0_15_ARCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_15_ARCACHE,
      twiddle_h_rsc_0_15_ARLOCK => twiddle_h_rsc_0_15_ARLOCK,
      twiddle_h_rsc_0_15_ARBURST => peaseNTT_core_inst_twiddle_h_rsc_0_15_ARBURST,
      twiddle_h_rsc_0_15_ARSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_15_ARSIZE,
      twiddle_h_rsc_0_15_ARLEN => peaseNTT_core_inst_twiddle_h_rsc_0_15_ARLEN,
      twiddle_h_rsc_0_15_ARADDR => peaseNTT_core_inst_twiddle_h_rsc_0_15_ARADDR,
      twiddle_h_rsc_0_15_ARID => twiddle_h_rsc_0_15_ARID,
      twiddle_h_rsc_0_15_BREADY => twiddle_h_rsc_0_15_BREADY,
      twiddle_h_rsc_0_15_BVALID => twiddle_h_rsc_0_15_BVALID,
      twiddle_h_rsc_0_15_BUSER => twiddle_h_rsc_0_15_BUSER,
      twiddle_h_rsc_0_15_BRESP => peaseNTT_core_inst_twiddle_h_rsc_0_15_BRESP,
      twiddle_h_rsc_0_15_BID => twiddle_h_rsc_0_15_BID,
      twiddle_h_rsc_0_15_WREADY => twiddle_h_rsc_0_15_WREADY,
      twiddle_h_rsc_0_15_WVALID => twiddle_h_rsc_0_15_WVALID,
      twiddle_h_rsc_0_15_WUSER => twiddle_h_rsc_0_15_WUSER,
      twiddle_h_rsc_0_15_WLAST => twiddle_h_rsc_0_15_WLAST,
      twiddle_h_rsc_0_15_WSTRB => peaseNTT_core_inst_twiddle_h_rsc_0_15_WSTRB,
      twiddle_h_rsc_0_15_WDATA => peaseNTT_core_inst_twiddle_h_rsc_0_15_WDATA,
      twiddle_h_rsc_0_15_AWREADY => twiddle_h_rsc_0_15_AWREADY,
      twiddle_h_rsc_0_15_AWVALID => twiddle_h_rsc_0_15_AWVALID,
      twiddle_h_rsc_0_15_AWUSER => twiddle_h_rsc_0_15_AWUSER,
      twiddle_h_rsc_0_15_AWREGION => peaseNTT_core_inst_twiddle_h_rsc_0_15_AWREGION,
      twiddle_h_rsc_0_15_AWQOS => peaseNTT_core_inst_twiddle_h_rsc_0_15_AWQOS,
      twiddle_h_rsc_0_15_AWPROT => peaseNTT_core_inst_twiddle_h_rsc_0_15_AWPROT,
      twiddle_h_rsc_0_15_AWCACHE => peaseNTT_core_inst_twiddle_h_rsc_0_15_AWCACHE,
      twiddle_h_rsc_0_15_AWLOCK => twiddle_h_rsc_0_15_AWLOCK,
      twiddle_h_rsc_0_15_AWBURST => peaseNTT_core_inst_twiddle_h_rsc_0_15_AWBURST,
      twiddle_h_rsc_0_15_AWSIZE => peaseNTT_core_inst_twiddle_h_rsc_0_15_AWSIZE,
      twiddle_h_rsc_0_15_AWLEN => peaseNTT_core_inst_twiddle_h_rsc_0_15_AWLEN,
      twiddle_h_rsc_0_15_AWADDR => peaseNTT_core_inst_twiddle_h_rsc_0_15_AWADDR,
      twiddle_h_rsc_0_15_AWID => twiddle_h_rsc_0_15_AWID,
      twiddle_h_rsc_triosy_0_15_lz => twiddle_h_rsc_triosy_0_15_lz,
      yt_rsc_0_0_i_clken_d => yt_rsc_0_0_i_clken_d,
      yt_rsc_0_0_i_qa_d => peaseNTT_core_inst_yt_rsc_0_0_i_qa_d,
      yt_rsc_0_1_i_qa_d => peaseNTT_core_inst_yt_rsc_0_1_i_qa_d,
      yt_rsc_0_2_i_qa_d => peaseNTT_core_inst_yt_rsc_0_2_i_qa_d,
      yt_rsc_0_3_i_qa_d => peaseNTT_core_inst_yt_rsc_0_3_i_qa_d,
      yt_rsc_0_4_i_qa_d => peaseNTT_core_inst_yt_rsc_0_4_i_qa_d,
      yt_rsc_0_5_i_qa_d => peaseNTT_core_inst_yt_rsc_0_5_i_qa_d,
      yt_rsc_0_6_i_qa_d => peaseNTT_core_inst_yt_rsc_0_6_i_qa_d,
      yt_rsc_0_7_i_qa_d => peaseNTT_core_inst_yt_rsc_0_7_i_qa_d,
      yt_rsc_0_8_i_qa_d => peaseNTT_core_inst_yt_rsc_0_8_i_qa_d,
      yt_rsc_0_9_i_qa_d => peaseNTT_core_inst_yt_rsc_0_9_i_qa_d,
      yt_rsc_0_10_i_qa_d => peaseNTT_core_inst_yt_rsc_0_10_i_qa_d,
      yt_rsc_0_11_i_qa_d => peaseNTT_core_inst_yt_rsc_0_11_i_qa_d,
      yt_rsc_0_12_i_qa_d => peaseNTT_core_inst_yt_rsc_0_12_i_qa_d,
      yt_rsc_0_13_i_qa_d => peaseNTT_core_inst_yt_rsc_0_13_i_qa_d,
      yt_rsc_0_14_i_qa_d => peaseNTT_core_inst_yt_rsc_0_14_i_qa_d,
      yt_rsc_0_15_i_qa_d => peaseNTT_core_inst_yt_rsc_0_15_i_qa_d,
      yt_rsc_0_16_i_clken_d => yt_rsc_0_16_i_clken_d,
      yt_rsc_0_16_i_qa_d => peaseNTT_core_inst_yt_rsc_0_16_i_qa_d,
      yt_rsc_0_17_i_qa_d => peaseNTT_core_inst_yt_rsc_0_17_i_qa_d,
      yt_rsc_0_18_i_qa_d => peaseNTT_core_inst_yt_rsc_0_18_i_qa_d,
      yt_rsc_0_19_i_qa_d => peaseNTT_core_inst_yt_rsc_0_19_i_qa_d,
      yt_rsc_0_20_i_qa_d => peaseNTT_core_inst_yt_rsc_0_20_i_qa_d,
      yt_rsc_0_21_i_qa_d => peaseNTT_core_inst_yt_rsc_0_21_i_qa_d,
      yt_rsc_0_22_i_qa_d => peaseNTT_core_inst_yt_rsc_0_22_i_qa_d,
      yt_rsc_0_23_i_qa_d => peaseNTT_core_inst_yt_rsc_0_23_i_qa_d,
      yt_rsc_0_24_i_qa_d => peaseNTT_core_inst_yt_rsc_0_24_i_qa_d,
      yt_rsc_0_25_i_qa_d => peaseNTT_core_inst_yt_rsc_0_25_i_qa_d,
      yt_rsc_0_26_i_qa_d => peaseNTT_core_inst_yt_rsc_0_26_i_qa_d,
      yt_rsc_0_27_i_qa_d => peaseNTT_core_inst_yt_rsc_0_27_i_qa_d,
      yt_rsc_0_28_i_qa_d => peaseNTT_core_inst_yt_rsc_0_28_i_qa_d,
      yt_rsc_0_29_i_qa_d => peaseNTT_core_inst_yt_rsc_0_29_i_qa_d,
      yt_rsc_0_30_i_qa_d => peaseNTT_core_inst_yt_rsc_0_30_i_qa_d,
      yt_rsc_0_31_i_qa_d => peaseNTT_core_inst_yt_rsc_0_31_i_qa_d,
      yt_rsc_1_0_i_clken_d => yt_rsc_1_0_i_clken_d,
      yt_rsc_1_0_i_da_d => peaseNTT_core_inst_yt_rsc_1_0_i_da_d,
      yt_rsc_1_0_i_qa_d => peaseNTT_core_inst_yt_rsc_1_0_i_qa_d,
      yt_rsc_1_1_i_da_d => peaseNTT_core_inst_yt_rsc_1_1_i_da_d,
      yt_rsc_1_1_i_qa_d => peaseNTT_core_inst_yt_rsc_1_1_i_qa_d,
      yt_rsc_1_2_i_da_d => peaseNTT_core_inst_yt_rsc_1_2_i_da_d,
      yt_rsc_1_2_i_qa_d => peaseNTT_core_inst_yt_rsc_1_2_i_qa_d,
      yt_rsc_1_3_i_da_d => peaseNTT_core_inst_yt_rsc_1_3_i_da_d,
      yt_rsc_1_3_i_qa_d => peaseNTT_core_inst_yt_rsc_1_3_i_qa_d,
      yt_rsc_1_4_i_da_d => peaseNTT_core_inst_yt_rsc_1_4_i_da_d,
      yt_rsc_1_4_i_qa_d => peaseNTT_core_inst_yt_rsc_1_4_i_qa_d,
      yt_rsc_1_5_i_da_d => peaseNTT_core_inst_yt_rsc_1_5_i_da_d,
      yt_rsc_1_5_i_qa_d => peaseNTT_core_inst_yt_rsc_1_5_i_qa_d,
      yt_rsc_1_6_i_da_d => peaseNTT_core_inst_yt_rsc_1_6_i_da_d,
      yt_rsc_1_6_i_qa_d => peaseNTT_core_inst_yt_rsc_1_6_i_qa_d,
      yt_rsc_1_7_i_da_d => peaseNTT_core_inst_yt_rsc_1_7_i_da_d,
      yt_rsc_1_7_i_qa_d => peaseNTT_core_inst_yt_rsc_1_7_i_qa_d,
      yt_rsc_1_8_i_da_d => peaseNTT_core_inst_yt_rsc_1_8_i_da_d,
      yt_rsc_1_8_i_qa_d => peaseNTT_core_inst_yt_rsc_1_8_i_qa_d,
      yt_rsc_1_9_i_da_d => peaseNTT_core_inst_yt_rsc_1_9_i_da_d,
      yt_rsc_1_9_i_qa_d => peaseNTT_core_inst_yt_rsc_1_9_i_qa_d,
      yt_rsc_1_10_i_da_d => peaseNTT_core_inst_yt_rsc_1_10_i_da_d,
      yt_rsc_1_10_i_qa_d => peaseNTT_core_inst_yt_rsc_1_10_i_qa_d,
      yt_rsc_1_11_i_da_d => peaseNTT_core_inst_yt_rsc_1_11_i_da_d,
      yt_rsc_1_11_i_qa_d => peaseNTT_core_inst_yt_rsc_1_11_i_qa_d,
      yt_rsc_1_12_i_da_d => peaseNTT_core_inst_yt_rsc_1_12_i_da_d,
      yt_rsc_1_12_i_qa_d => peaseNTT_core_inst_yt_rsc_1_12_i_qa_d,
      yt_rsc_1_13_i_da_d => peaseNTT_core_inst_yt_rsc_1_13_i_da_d,
      yt_rsc_1_13_i_qa_d => peaseNTT_core_inst_yt_rsc_1_13_i_qa_d,
      yt_rsc_1_14_i_da_d => peaseNTT_core_inst_yt_rsc_1_14_i_da_d,
      yt_rsc_1_14_i_qa_d => peaseNTT_core_inst_yt_rsc_1_14_i_qa_d,
      yt_rsc_1_15_i_da_d => peaseNTT_core_inst_yt_rsc_1_15_i_da_d,
      yt_rsc_1_15_i_qa_d => peaseNTT_core_inst_yt_rsc_1_15_i_qa_d,
      yt_rsc_1_16_i_clken_d => yt_rsc_1_16_i_clken_d,
      yt_rsc_1_16_i_da_d => peaseNTT_core_inst_yt_rsc_1_16_i_da_d,
      yt_rsc_1_16_i_qa_d => peaseNTT_core_inst_yt_rsc_1_16_i_qa_d,
      yt_rsc_1_17_i_da_d => peaseNTT_core_inst_yt_rsc_1_17_i_da_d,
      yt_rsc_1_17_i_qa_d => peaseNTT_core_inst_yt_rsc_1_17_i_qa_d,
      yt_rsc_1_18_i_da_d => peaseNTT_core_inst_yt_rsc_1_18_i_da_d,
      yt_rsc_1_18_i_qa_d => peaseNTT_core_inst_yt_rsc_1_18_i_qa_d,
      yt_rsc_1_19_i_da_d => peaseNTT_core_inst_yt_rsc_1_19_i_da_d,
      yt_rsc_1_19_i_qa_d => peaseNTT_core_inst_yt_rsc_1_19_i_qa_d,
      yt_rsc_1_20_i_da_d => peaseNTT_core_inst_yt_rsc_1_20_i_da_d,
      yt_rsc_1_20_i_qa_d => peaseNTT_core_inst_yt_rsc_1_20_i_qa_d,
      yt_rsc_1_21_i_da_d => peaseNTT_core_inst_yt_rsc_1_21_i_da_d,
      yt_rsc_1_21_i_qa_d => peaseNTT_core_inst_yt_rsc_1_21_i_qa_d,
      yt_rsc_1_22_i_da_d => peaseNTT_core_inst_yt_rsc_1_22_i_da_d,
      yt_rsc_1_22_i_qa_d => peaseNTT_core_inst_yt_rsc_1_22_i_qa_d,
      yt_rsc_1_23_i_da_d => peaseNTT_core_inst_yt_rsc_1_23_i_da_d,
      yt_rsc_1_23_i_qa_d => peaseNTT_core_inst_yt_rsc_1_23_i_qa_d,
      yt_rsc_1_24_i_da_d => peaseNTT_core_inst_yt_rsc_1_24_i_da_d,
      yt_rsc_1_24_i_qa_d => peaseNTT_core_inst_yt_rsc_1_24_i_qa_d,
      yt_rsc_1_25_i_da_d => peaseNTT_core_inst_yt_rsc_1_25_i_da_d,
      yt_rsc_1_25_i_qa_d => peaseNTT_core_inst_yt_rsc_1_25_i_qa_d,
      yt_rsc_1_26_i_da_d => peaseNTT_core_inst_yt_rsc_1_26_i_da_d,
      yt_rsc_1_26_i_qa_d => peaseNTT_core_inst_yt_rsc_1_26_i_qa_d,
      yt_rsc_1_27_i_da_d => peaseNTT_core_inst_yt_rsc_1_27_i_da_d,
      yt_rsc_1_27_i_qa_d => peaseNTT_core_inst_yt_rsc_1_27_i_qa_d,
      yt_rsc_1_28_i_da_d => peaseNTT_core_inst_yt_rsc_1_28_i_da_d,
      yt_rsc_1_28_i_qa_d => peaseNTT_core_inst_yt_rsc_1_28_i_qa_d,
      yt_rsc_1_29_i_da_d => peaseNTT_core_inst_yt_rsc_1_29_i_da_d,
      yt_rsc_1_29_i_qa_d => peaseNTT_core_inst_yt_rsc_1_29_i_qa_d,
      yt_rsc_1_30_i_da_d => peaseNTT_core_inst_yt_rsc_1_30_i_da_d,
      yt_rsc_1_30_i_qa_d => peaseNTT_core_inst_yt_rsc_1_30_i_qa_d,
      yt_rsc_1_31_i_da_d => peaseNTT_core_inst_yt_rsc_1_31_i_da_d,
      yt_rsc_1_31_i_qa_d => peaseNTT_core_inst_yt_rsc_1_31_i_qa_d,
      xt_rsc_0_0_i_qa_d => peaseNTT_core_inst_xt_rsc_0_0_i_qa_d,
      xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_1_i_qa_d => peaseNTT_core_inst_xt_rsc_0_1_i_qa_d,
      xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_2_i_qa_d => peaseNTT_core_inst_xt_rsc_0_2_i_qa_d,
      xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_3_i_qa_d => peaseNTT_core_inst_xt_rsc_0_3_i_qa_d,
      xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_4_i_qa_d => peaseNTT_core_inst_xt_rsc_0_4_i_qa_d,
      xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_5_i_qa_d => peaseNTT_core_inst_xt_rsc_0_5_i_qa_d,
      xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_6_i_qa_d => peaseNTT_core_inst_xt_rsc_0_6_i_qa_d,
      xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_7_i_qa_d => peaseNTT_core_inst_xt_rsc_0_7_i_qa_d,
      xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_8_i_qa_d => peaseNTT_core_inst_xt_rsc_0_8_i_qa_d,
      xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_9_i_qa_d => peaseNTT_core_inst_xt_rsc_0_9_i_qa_d,
      xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_10_i_qa_d => peaseNTT_core_inst_xt_rsc_0_10_i_qa_d,
      xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_11_i_qa_d => peaseNTT_core_inst_xt_rsc_0_11_i_qa_d,
      xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_12_i_qa_d => peaseNTT_core_inst_xt_rsc_0_12_i_qa_d,
      xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_13_i_qa_d => peaseNTT_core_inst_xt_rsc_0_13_i_qa_d,
      xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_14_i_qa_d => peaseNTT_core_inst_xt_rsc_0_14_i_qa_d,
      xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_15_i_qa_d => peaseNTT_core_inst_xt_rsc_0_15_i_qa_d,
      xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_16_i_qa_d => peaseNTT_core_inst_xt_rsc_0_16_i_qa_d,
      xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_16_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_17_i_qa_d => peaseNTT_core_inst_xt_rsc_0_17_i_qa_d,
      xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_17_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_18_i_qa_d => peaseNTT_core_inst_xt_rsc_0_18_i_qa_d,
      xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_18_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_19_i_qa_d => peaseNTT_core_inst_xt_rsc_0_19_i_qa_d,
      xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_19_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_20_i_qa_d => peaseNTT_core_inst_xt_rsc_0_20_i_qa_d,
      xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_20_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_21_i_qa_d => peaseNTT_core_inst_xt_rsc_0_21_i_qa_d,
      xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_21_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_22_i_qa_d => peaseNTT_core_inst_xt_rsc_0_22_i_qa_d,
      xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_22_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_23_i_qa_d => peaseNTT_core_inst_xt_rsc_0_23_i_qa_d,
      xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_23_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_24_i_qa_d => peaseNTT_core_inst_xt_rsc_0_24_i_qa_d,
      xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_24_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_25_i_qa_d => peaseNTT_core_inst_xt_rsc_0_25_i_qa_d,
      xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_25_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_26_i_qa_d => peaseNTT_core_inst_xt_rsc_0_26_i_qa_d,
      xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_26_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_27_i_qa_d => peaseNTT_core_inst_xt_rsc_0_27_i_qa_d,
      xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_27_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_28_i_qa_d => peaseNTT_core_inst_xt_rsc_0_28_i_qa_d,
      xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_28_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_29_i_qa_d => peaseNTT_core_inst_xt_rsc_0_29_i_qa_d,
      xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_29_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_30_i_qa_d => peaseNTT_core_inst_xt_rsc_0_30_i_qa_d,
      xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_30_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_0_31_i_qa_d => peaseNTT_core_inst_xt_rsc_0_31_i_qa_d,
      xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_0_31_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_0_i_qa_d => peaseNTT_core_inst_xt_rsc_1_0_i_qa_d,
      xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_1_i_qa_d => peaseNTT_core_inst_xt_rsc_1_1_i_qa_d,
      xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_1_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_2_i_qa_d => peaseNTT_core_inst_xt_rsc_1_2_i_qa_d,
      xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_2_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_3_i_qa_d => peaseNTT_core_inst_xt_rsc_1_3_i_qa_d,
      xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_3_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_4_i_qa_d => peaseNTT_core_inst_xt_rsc_1_4_i_qa_d,
      xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_4_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_5_i_qa_d => peaseNTT_core_inst_xt_rsc_1_5_i_qa_d,
      xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_5_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_6_i_qa_d => peaseNTT_core_inst_xt_rsc_1_6_i_qa_d,
      xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_6_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_7_i_qa_d => peaseNTT_core_inst_xt_rsc_1_7_i_qa_d,
      xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_7_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_8_i_qa_d => peaseNTT_core_inst_xt_rsc_1_8_i_qa_d,
      xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_8_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_9_i_qa_d => peaseNTT_core_inst_xt_rsc_1_9_i_qa_d,
      xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_9_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_10_i_qa_d => peaseNTT_core_inst_xt_rsc_1_10_i_qa_d,
      xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_10_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_11_i_qa_d => peaseNTT_core_inst_xt_rsc_1_11_i_qa_d,
      xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_11_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_12_i_qa_d => peaseNTT_core_inst_xt_rsc_1_12_i_qa_d,
      xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_12_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_13_i_qa_d => peaseNTT_core_inst_xt_rsc_1_13_i_qa_d,
      xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_13_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_14_i_qa_d => peaseNTT_core_inst_xt_rsc_1_14_i_qa_d,
      xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_14_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_15_i_qa_d => peaseNTT_core_inst_xt_rsc_1_15_i_qa_d,
      xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_15_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_16_i_qa_d => peaseNTT_core_inst_xt_rsc_1_16_i_qa_d,
      xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_16_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_17_i_qa_d => peaseNTT_core_inst_xt_rsc_1_17_i_qa_d,
      xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_17_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_18_i_qa_d => peaseNTT_core_inst_xt_rsc_1_18_i_qa_d,
      xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_18_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_19_i_qa_d => peaseNTT_core_inst_xt_rsc_1_19_i_qa_d,
      xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_19_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_20_i_qa_d => peaseNTT_core_inst_xt_rsc_1_20_i_qa_d,
      xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_20_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_21_i_qa_d => peaseNTT_core_inst_xt_rsc_1_21_i_qa_d,
      xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_21_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_22_i_qa_d => peaseNTT_core_inst_xt_rsc_1_22_i_qa_d,
      xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_22_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_23_i_qa_d => peaseNTT_core_inst_xt_rsc_1_23_i_qa_d,
      xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_23_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_24_i_qa_d => peaseNTT_core_inst_xt_rsc_1_24_i_qa_d,
      xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_24_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_25_i_qa_d => peaseNTT_core_inst_xt_rsc_1_25_i_qa_d,
      xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_25_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_26_i_qa_d => peaseNTT_core_inst_xt_rsc_1_26_i_qa_d,
      xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_26_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_27_i_qa_d => peaseNTT_core_inst_xt_rsc_1_27_i_qa_d,
      xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_27_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_28_i_qa_d => peaseNTT_core_inst_xt_rsc_1_28_i_qa_d,
      xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_28_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_29_i_qa_d => peaseNTT_core_inst_xt_rsc_1_29_i_qa_d,
      xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_29_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_30_i_qa_d => peaseNTT_core_inst_xt_rsc_1_30_i_qa_d,
      xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_30_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      xt_rsc_1_31_i_qa_d => peaseNTT_core_inst_xt_rsc_1_31_i_qa_d,
      xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d => xt_rsc_1_31_i_rwA_rw_ram_ir_internal_RMASK_B_d,
      yt_rsc_0_0_i_adra_d_pff => peaseNTT_core_inst_yt_rsc_0_0_i_adra_d_pff,
      yt_rsc_0_0_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_0_i_da_d_pff,
      yt_rsc_0_0_i_wea_d_pff => yt_rsc_0_0_i_wea_d_iff,
      yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff => yt_rsc_0_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      yt_rsc_0_1_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_1_i_da_d_pff,
      yt_rsc_0_2_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_2_i_da_d_pff,
      yt_rsc_0_3_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_3_i_da_d_pff,
      yt_rsc_0_4_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_4_i_da_d_pff,
      yt_rsc_0_5_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_5_i_da_d_pff,
      yt_rsc_0_6_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_6_i_da_d_pff,
      yt_rsc_0_7_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_7_i_da_d_pff,
      yt_rsc_0_8_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_8_i_da_d_pff,
      yt_rsc_0_9_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_9_i_da_d_pff,
      yt_rsc_0_10_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_10_i_da_d_pff,
      yt_rsc_0_11_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_11_i_da_d_pff,
      yt_rsc_0_12_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_12_i_da_d_pff,
      yt_rsc_0_13_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_13_i_da_d_pff,
      yt_rsc_0_14_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_14_i_da_d_pff,
      yt_rsc_0_15_i_da_d_pff => peaseNTT_core_inst_yt_rsc_0_15_i_da_d_pff,
      yt_rsc_0_16_i_adra_d_pff => peaseNTT_core_inst_yt_rsc_0_16_i_adra_d_pff,
      yt_rsc_0_16_i_wea_d_pff => yt_rsc_0_16_i_wea_d_iff,
      yt_rsc_1_0_i_adra_d_pff => peaseNTT_core_inst_yt_rsc_1_0_i_adra_d_pff,
      yt_rsc_1_0_i_wea_d_pff => yt_rsc_1_0_i_wea_d_iff,
      yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_pff => yt_rsc_1_0_i_rwA_rw_ram_ir_internal_RMASK_B_d_iff,
      yt_rsc_1_16_i_adra_d_pff => peaseNTT_core_inst_yt_rsc_1_16_i_adra_d_pff,
      yt_rsc_1_16_i_wea_d_pff => yt_rsc_1_16_i_wea_d_iff,
      xt_rsc_0_0_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_0_i_adra_d_pff,
      xt_rsc_0_0_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_0_i_da_d_pff,
      xt_rsc_0_0_i_wea_d_pff => xt_rsc_0_0_i_wea_d_iff,
      xt_rsc_0_1_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_1_i_da_d_pff,
      xt_rsc_0_1_i_wea_d_pff => xt_rsc_0_1_i_wea_d_iff,
      xt_rsc_0_2_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_2_i_da_d_pff,
      xt_rsc_0_2_i_wea_d_pff => xt_rsc_0_2_i_wea_d_iff,
      xt_rsc_0_3_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_3_i_da_d_pff,
      xt_rsc_0_3_i_wea_d_pff => xt_rsc_0_3_i_wea_d_iff,
      xt_rsc_0_4_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_4_i_da_d_pff,
      xt_rsc_0_4_i_wea_d_pff => xt_rsc_0_4_i_wea_d_iff,
      xt_rsc_0_5_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_5_i_da_d_pff,
      xt_rsc_0_5_i_wea_d_pff => xt_rsc_0_5_i_wea_d_iff,
      xt_rsc_0_6_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_6_i_da_d_pff,
      xt_rsc_0_6_i_wea_d_pff => xt_rsc_0_6_i_wea_d_iff,
      xt_rsc_0_7_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_7_i_da_d_pff,
      xt_rsc_0_7_i_wea_d_pff => xt_rsc_0_7_i_wea_d_iff,
      xt_rsc_0_8_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_8_i_da_d_pff,
      xt_rsc_0_8_i_wea_d_pff => xt_rsc_0_8_i_wea_d_iff,
      xt_rsc_0_9_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_9_i_da_d_pff,
      xt_rsc_0_9_i_wea_d_pff => xt_rsc_0_9_i_wea_d_iff,
      xt_rsc_0_10_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_10_i_da_d_pff,
      xt_rsc_0_10_i_wea_d_pff => xt_rsc_0_10_i_wea_d_iff,
      xt_rsc_0_11_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_11_i_da_d_pff,
      xt_rsc_0_11_i_wea_d_pff => xt_rsc_0_11_i_wea_d_iff,
      xt_rsc_0_12_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_12_i_da_d_pff,
      xt_rsc_0_12_i_wea_d_pff => xt_rsc_0_12_i_wea_d_iff,
      xt_rsc_0_13_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_13_i_da_d_pff,
      xt_rsc_0_13_i_wea_d_pff => xt_rsc_0_13_i_wea_d_iff,
      xt_rsc_0_14_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_14_i_da_d_pff,
      xt_rsc_0_14_i_wea_d_pff => xt_rsc_0_14_i_wea_d_iff,
      xt_rsc_0_15_i_da_d_pff => peaseNTT_core_inst_xt_rsc_0_15_i_da_d_pff,
      xt_rsc_0_15_i_wea_d_pff => xt_rsc_0_15_i_wea_d_iff,
      xt_rsc_0_16_i_adra_d_pff => peaseNTT_core_inst_xt_rsc_0_16_i_adra_d_pff,
      xt_rsc_0_16_i_wea_d_pff => xt_rsc_0_16_i_wea_d_iff,
      xt_rsc_0_17_i_wea_d_pff => xt_rsc_0_17_i_wea_d_iff,
      xt_rsc_0_18_i_wea_d_pff => xt_rsc_0_18_i_wea_d_iff,
      xt_rsc_0_19_i_wea_d_pff => xt_rsc_0_19_i_wea_d_iff,
      xt_rsc_0_20_i_wea_d_pff => xt_rsc_0_20_i_wea_d_iff,
      xt_rsc_0_21_i_wea_d_pff => xt_rsc_0_21_i_wea_d_iff,
      xt_rsc_0_22_i_wea_d_pff => xt_rsc_0_22_i_wea_d_iff,
      xt_rsc_0_23_i_wea_d_pff => xt_rsc_0_23_i_wea_d_iff,
      xt_rsc_0_24_i_wea_d_pff => xt_rsc_0_24_i_wea_d_iff,
      xt_rsc_0_25_i_wea_d_pff => xt_rsc_0_25_i_wea_d_iff,
      xt_rsc_0_26_i_wea_d_pff => xt_rsc_0_26_i_wea_d_iff,
      xt_rsc_0_27_i_wea_d_pff => xt_rsc_0_27_i_wea_d_iff,
      xt_rsc_0_28_i_wea_d_pff => xt_rsc_0_28_i_wea_d_iff,
      xt_rsc_0_29_i_wea_d_pff => xt_rsc_0_29_i_wea_d_iff,
      xt_rsc_0_30_i_wea_d_pff => xt_rsc_0_30_i_wea_d_iff,
      xt_rsc_0_31_i_wea_d_pff => xt_rsc_0_31_i_wea_d_iff,
      xt_rsc_1_0_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_0_i_da_d_pff,
      xt_rsc_1_0_i_wea_d_pff => xt_rsc_1_0_i_wea_d_iff,
      xt_rsc_1_1_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_1_i_da_d_pff,
      xt_rsc_1_1_i_wea_d_pff => xt_rsc_1_1_i_wea_d_iff,
      xt_rsc_1_2_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_2_i_da_d_pff,
      xt_rsc_1_2_i_wea_d_pff => xt_rsc_1_2_i_wea_d_iff,
      xt_rsc_1_3_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_3_i_da_d_pff,
      xt_rsc_1_3_i_wea_d_pff => xt_rsc_1_3_i_wea_d_iff,
      xt_rsc_1_4_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_4_i_da_d_pff,
      xt_rsc_1_4_i_wea_d_pff => xt_rsc_1_4_i_wea_d_iff,
      xt_rsc_1_5_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_5_i_da_d_pff,
      xt_rsc_1_5_i_wea_d_pff => xt_rsc_1_5_i_wea_d_iff,
      xt_rsc_1_6_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_6_i_da_d_pff,
      xt_rsc_1_6_i_wea_d_pff => xt_rsc_1_6_i_wea_d_iff,
      xt_rsc_1_7_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_7_i_da_d_pff,
      xt_rsc_1_7_i_wea_d_pff => xt_rsc_1_7_i_wea_d_iff,
      xt_rsc_1_8_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_8_i_da_d_pff,
      xt_rsc_1_8_i_wea_d_pff => xt_rsc_1_8_i_wea_d_iff,
      xt_rsc_1_9_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_9_i_da_d_pff,
      xt_rsc_1_9_i_wea_d_pff => xt_rsc_1_9_i_wea_d_iff,
      xt_rsc_1_10_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_10_i_da_d_pff,
      xt_rsc_1_10_i_wea_d_pff => xt_rsc_1_10_i_wea_d_iff,
      xt_rsc_1_11_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_11_i_da_d_pff,
      xt_rsc_1_11_i_wea_d_pff => xt_rsc_1_11_i_wea_d_iff,
      xt_rsc_1_12_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_12_i_da_d_pff,
      xt_rsc_1_12_i_wea_d_pff => xt_rsc_1_12_i_wea_d_iff,
      xt_rsc_1_13_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_13_i_da_d_pff,
      xt_rsc_1_13_i_wea_d_pff => xt_rsc_1_13_i_wea_d_iff,
      xt_rsc_1_14_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_14_i_da_d_pff,
      xt_rsc_1_14_i_wea_d_pff => xt_rsc_1_14_i_wea_d_iff,
      xt_rsc_1_15_i_da_d_pff => peaseNTT_core_inst_xt_rsc_1_15_i_da_d_pff,
      xt_rsc_1_15_i_wea_d_pff => xt_rsc_1_15_i_wea_d_iff,
      xt_rsc_1_16_i_wea_d_pff => xt_rsc_1_16_i_wea_d_iff,
      xt_rsc_1_17_i_wea_d_pff => xt_rsc_1_17_i_wea_d_iff,
      xt_rsc_1_18_i_wea_d_pff => xt_rsc_1_18_i_wea_d_iff,
      xt_rsc_1_19_i_wea_d_pff => xt_rsc_1_19_i_wea_d_iff,
      xt_rsc_1_20_i_wea_d_pff => xt_rsc_1_20_i_wea_d_iff,
      xt_rsc_1_21_i_wea_d_pff => xt_rsc_1_21_i_wea_d_iff,
      xt_rsc_1_22_i_wea_d_pff => xt_rsc_1_22_i_wea_d_iff,
      xt_rsc_1_23_i_wea_d_pff => xt_rsc_1_23_i_wea_d_iff,
      xt_rsc_1_24_i_wea_d_pff => xt_rsc_1_24_i_wea_d_iff,
      xt_rsc_1_25_i_wea_d_pff => xt_rsc_1_25_i_wea_d_iff,
      xt_rsc_1_26_i_wea_d_pff => xt_rsc_1_26_i_wea_d_iff,
      xt_rsc_1_27_i_wea_d_pff => xt_rsc_1_27_i_wea_d_iff,
      xt_rsc_1_28_i_wea_d_pff => xt_rsc_1_28_i_wea_d_iff,
      xt_rsc_1_29_i_wea_d_pff => xt_rsc_1_29_i_wea_d_iff,
      xt_rsc_1_30_i_wea_d_pff => xt_rsc_1_30_i_wea_d_iff,
      xt_rsc_1_31_i_wea_d_pff => xt_rsc_1_31_i_wea_d_iff
    );
  peaseNTT_core_inst_p_rsc_dat <= p_rsc_dat;
  twiddle_rsc_0_0_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_0_RRESP;
  twiddle_rsc_0_0_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_0_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_0_ARREGION <= twiddle_rsc_0_0_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_0_ARQOS <= twiddle_rsc_0_0_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_0_ARPROT <= twiddle_rsc_0_0_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_0_ARCACHE <= twiddle_rsc_0_0_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_0_ARBURST <= twiddle_rsc_0_0_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_0_ARSIZE <= twiddle_rsc_0_0_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_0_ARLEN <= twiddle_rsc_0_0_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_0_ARADDR <= twiddle_rsc_0_0_ARADDR;
  twiddle_rsc_0_0_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_0_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_0_WSTRB <= twiddle_rsc_0_0_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_0_WDATA <= twiddle_rsc_0_0_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_0_AWREGION <= twiddle_rsc_0_0_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_0_AWQOS <= twiddle_rsc_0_0_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_0_AWPROT <= twiddle_rsc_0_0_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_0_AWCACHE <= twiddle_rsc_0_0_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_0_AWBURST <= twiddle_rsc_0_0_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_0_AWSIZE <= twiddle_rsc_0_0_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_0_AWLEN <= twiddle_rsc_0_0_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_0_AWADDR <= twiddle_rsc_0_0_AWADDR;
  twiddle_rsc_0_1_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_1_RRESP;
  twiddle_rsc_0_1_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_1_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_1_ARREGION <= twiddle_rsc_0_1_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_1_ARQOS <= twiddle_rsc_0_1_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_1_ARPROT <= twiddle_rsc_0_1_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_1_ARCACHE <= twiddle_rsc_0_1_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_1_ARBURST <= twiddle_rsc_0_1_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_1_ARSIZE <= twiddle_rsc_0_1_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_1_ARLEN <= twiddle_rsc_0_1_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_1_ARADDR <= twiddle_rsc_0_1_ARADDR;
  twiddle_rsc_0_1_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_1_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_1_WSTRB <= twiddle_rsc_0_1_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_1_WDATA <= twiddle_rsc_0_1_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_1_AWREGION <= twiddle_rsc_0_1_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_1_AWQOS <= twiddle_rsc_0_1_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_1_AWPROT <= twiddle_rsc_0_1_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_1_AWCACHE <= twiddle_rsc_0_1_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_1_AWBURST <= twiddle_rsc_0_1_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_1_AWSIZE <= twiddle_rsc_0_1_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_1_AWLEN <= twiddle_rsc_0_1_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_1_AWADDR <= twiddle_rsc_0_1_AWADDR;
  twiddle_rsc_0_2_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_2_RRESP;
  twiddle_rsc_0_2_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_2_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_2_ARREGION <= twiddle_rsc_0_2_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_2_ARQOS <= twiddle_rsc_0_2_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_2_ARPROT <= twiddle_rsc_0_2_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_2_ARCACHE <= twiddle_rsc_0_2_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_2_ARBURST <= twiddle_rsc_0_2_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_2_ARSIZE <= twiddle_rsc_0_2_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_2_ARLEN <= twiddle_rsc_0_2_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_2_ARADDR <= twiddle_rsc_0_2_ARADDR;
  twiddle_rsc_0_2_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_2_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_2_WSTRB <= twiddle_rsc_0_2_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_2_WDATA <= twiddle_rsc_0_2_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_2_AWREGION <= twiddle_rsc_0_2_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_2_AWQOS <= twiddle_rsc_0_2_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_2_AWPROT <= twiddle_rsc_0_2_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_2_AWCACHE <= twiddle_rsc_0_2_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_2_AWBURST <= twiddle_rsc_0_2_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_2_AWSIZE <= twiddle_rsc_0_2_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_2_AWLEN <= twiddle_rsc_0_2_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_2_AWADDR <= twiddle_rsc_0_2_AWADDR;
  twiddle_rsc_0_3_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_3_RRESP;
  twiddle_rsc_0_3_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_3_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_3_ARREGION <= twiddle_rsc_0_3_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_3_ARQOS <= twiddle_rsc_0_3_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_3_ARPROT <= twiddle_rsc_0_3_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_3_ARCACHE <= twiddle_rsc_0_3_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_3_ARBURST <= twiddle_rsc_0_3_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_3_ARSIZE <= twiddle_rsc_0_3_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_3_ARLEN <= twiddle_rsc_0_3_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_3_ARADDR <= twiddle_rsc_0_3_ARADDR;
  twiddle_rsc_0_3_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_3_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_3_WSTRB <= twiddle_rsc_0_3_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_3_WDATA <= twiddle_rsc_0_3_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_3_AWREGION <= twiddle_rsc_0_3_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_3_AWQOS <= twiddle_rsc_0_3_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_3_AWPROT <= twiddle_rsc_0_3_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_3_AWCACHE <= twiddle_rsc_0_3_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_3_AWBURST <= twiddle_rsc_0_3_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_3_AWSIZE <= twiddle_rsc_0_3_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_3_AWLEN <= twiddle_rsc_0_3_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_3_AWADDR <= twiddle_rsc_0_3_AWADDR;
  twiddle_rsc_0_4_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_4_RRESP;
  twiddle_rsc_0_4_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_4_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_4_ARREGION <= twiddle_rsc_0_4_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_4_ARQOS <= twiddle_rsc_0_4_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_4_ARPROT <= twiddle_rsc_0_4_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_4_ARCACHE <= twiddle_rsc_0_4_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_4_ARBURST <= twiddle_rsc_0_4_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_4_ARSIZE <= twiddle_rsc_0_4_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_4_ARLEN <= twiddle_rsc_0_4_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_4_ARADDR <= twiddle_rsc_0_4_ARADDR;
  twiddle_rsc_0_4_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_4_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_4_WSTRB <= twiddle_rsc_0_4_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_4_WDATA <= twiddle_rsc_0_4_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_4_AWREGION <= twiddle_rsc_0_4_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_4_AWQOS <= twiddle_rsc_0_4_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_4_AWPROT <= twiddle_rsc_0_4_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_4_AWCACHE <= twiddle_rsc_0_4_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_4_AWBURST <= twiddle_rsc_0_4_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_4_AWSIZE <= twiddle_rsc_0_4_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_4_AWLEN <= twiddle_rsc_0_4_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_4_AWADDR <= twiddle_rsc_0_4_AWADDR;
  twiddle_rsc_0_5_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_5_RRESP;
  twiddle_rsc_0_5_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_5_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_5_ARREGION <= twiddle_rsc_0_5_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_5_ARQOS <= twiddle_rsc_0_5_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_5_ARPROT <= twiddle_rsc_0_5_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_5_ARCACHE <= twiddle_rsc_0_5_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_5_ARBURST <= twiddle_rsc_0_5_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_5_ARSIZE <= twiddle_rsc_0_5_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_5_ARLEN <= twiddle_rsc_0_5_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_5_ARADDR <= twiddle_rsc_0_5_ARADDR;
  twiddle_rsc_0_5_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_5_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_5_WSTRB <= twiddle_rsc_0_5_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_5_WDATA <= twiddle_rsc_0_5_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_5_AWREGION <= twiddle_rsc_0_5_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_5_AWQOS <= twiddle_rsc_0_5_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_5_AWPROT <= twiddle_rsc_0_5_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_5_AWCACHE <= twiddle_rsc_0_5_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_5_AWBURST <= twiddle_rsc_0_5_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_5_AWSIZE <= twiddle_rsc_0_5_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_5_AWLEN <= twiddle_rsc_0_5_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_5_AWADDR <= twiddle_rsc_0_5_AWADDR;
  twiddle_rsc_0_6_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_6_RRESP;
  twiddle_rsc_0_6_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_6_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_6_ARREGION <= twiddle_rsc_0_6_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_6_ARQOS <= twiddle_rsc_0_6_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_6_ARPROT <= twiddle_rsc_0_6_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_6_ARCACHE <= twiddle_rsc_0_6_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_6_ARBURST <= twiddle_rsc_0_6_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_6_ARSIZE <= twiddle_rsc_0_6_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_6_ARLEN <= twiddle_rsc_0_6_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_6_ARADDR <= twiddle_rsc_0_6_ARADDR;
  twiddle_rsc_0_6_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_6_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_6_WSTRB <= twiddle_rsc_0_6_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_6_WDATA <= twiddle_rsc_0_6_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_6_AWREGION <= twiddle_rsc_0_6_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_6_AWQOS <= twiddle_rsc_0_6_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_6_AWPROT <= twiddle_rsc_0_6_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_6_AWCACHE <= twiddle_rsc_0_6_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_6_AWBURST <= twiddle_rsc_0_6_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_6_AWSIZE <= twiddle_rsc_0_6_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_6_AWLEN <= twiddle_rsc_0_6_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_6_AWADDR <= twiddle_rsc_0_6_AWADDR;
  twiddle_rsc_0_7_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_7_RRESP;
  twiddle_rsc_0_7_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_7_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_7_ARREGION <= twiddle_rsc_0_7_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_7_ARQOS <= twiddle_rsc_0_7_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_7_ARPROT <= twiddle_rsc_0_7_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_7_ARCACHE <= twiddle_rsc_0_7_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_7_ARBURST <= twiddle_rsc_0_7_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_7_ARSIZE <= twiddle_rsc_0_7_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_7_ARLEN <= twiddle_rsc_0_7_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_7_ARADDR <= twiddle_rsc_0_7_ARADDR;
  twiddle_rsc_0_7_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_7_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_7_WSTRB <= twiddle_rsc_0_7_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_7_WDATA <= twiddle_rsc_0_7_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_7_AWREGION <= twiddle_rsc_0_7_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_7_AWQOS <= twiddle_rsc_0_7_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_7_AWPROT <= twiddle_rsc_0_7_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_7_AWCACHE <= twiddle_rsc_0_7_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_7_AWBURST <= twiddle_rsc_0_7_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_7_AWSIZE <= twiddle_rsc_0_7_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_7_AWLEN <= twiddle_rsc_0_7_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_7_AWADDR <= twiddle_rsc_0_7_AWADDR;
  twiddle_rsc_0_8_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_8_RRESP;
  twiddle_rsc_0_8_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_8_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_8_ARREGION <= twiddle_rsc_0_8_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_8_ARQOS <= twiddle_rsc_0_8_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_8_ARPROT <= twiddle_rsc_0_8_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_8_ARCACHE <= twiddle_rsc_0_8_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_8_ARBURST <= twiddle_rsc_0_8_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_8_ARSIZE <= twiddle_rsc_0_8_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_8_ARLEN <= twiddle_rsc_0_8_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_8_ARADDR <= twiddle_rsc_0_8_ARADDR;
  twiddle_rsc_0_8_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_8_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_8_WSTRB <= twiddle_rsc_0_8_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_8_WDATA <= twiddle_rsc_0_8_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_8_AWREGION <= twiddle_rsc_0_8_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_8_AWQOS <= twiddle_rsc_0_8_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_8_AWPROT <= twiddle_rsc_0_8_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_8_AWCACHE <= twiddle_rsc_0_8_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_8_AWBURST <= twiddle_rsc_0_8_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_8_AWSIZE <= twiddle_rsc_0_8_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_8_AWLEN <= twiddle_rsc_0_8_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_8_AWADDR <= twiddle_rsc_0_8_AWADDR;
  twiddle_rsc_0_9_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_9_RRESP;
  twiddle_rsc_0_9_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_9_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_9_ARREGION <= twiddle_rsc_0_9_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_9_ARQOS <= twiddle_rsc_0_9_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_9_ARPROT <= twiddle_rsc_0_9_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_9_ARCACHE <= twiddle_rsc_0_9_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_9_ARBURST <= twiddle_rsc_0_9_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_9_ARSIZE <= twiddle_rsc_0_9_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_9_ARLEN <= twiddle_rsc_0_9_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_9_ARADDR <= twiddle_rsc_0_9_ARADDR;
  twiddle_rsc_0_9_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_9_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_9_WSTRB <= twiddle_rsc_0_9_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_9_WDATA <= twiddle_rsc_0_9_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_9_AWREGION <= twiddle_rsc_0_9_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_9_AWQOS <= twiddle_rsc_0_9_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_9_AWPROT <= twiddle_rsc_0_9_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_9_AWCACHE <= twiddle_rsc_0_9_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_9_AWBURST <= twiddle_rsc_0_9_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_9_AWSIZE <= twiddle_rsc_0_9_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_9_AWLEN <= twiddle_rsc_0_9_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_9_AWADDR <= twiddle_rsc_0_9_AWADDR;
  twiddle_rsc_0_10_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_10_RRESP;
  twiddle_rsc_0_10_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_10_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_10_ARREGION <= twiddle_rsc_0_10_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_10_ARQOS <= twiddle_rsc_0_10_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_10_ARPROT <= twiddle_rsc_0_10_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_10_ARCACHE <= twiddle_rsc_0_10_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_10_ARBURST <= twiddle_rsc_0_10_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_10_ARSIZE <= twiddle_rsc_0_10_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_10_ARLEN <= twiddle_rsc_0_10_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_10_ARADDR <= twiddle_rsc_0_10_ARADDR;
  twiddle_rsc_0_10_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_10_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_10_WSTRB <= twiddle_rsc_0_10_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_10_WDATA <= twiddle_rsc_0_10_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_10_AWREGION <= twiddle_rsc_0_10_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_10_AWQOS <= twiddle_rsc_0_10_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_10_AWPROT <= twiddle_rsc_0_10_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_10_AWCACHE <= twiddle_rsc_0_10_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_10_AWBURST <= twiddle_rsc_0_10_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_10_AWSIZE <= twiddle_rsc_0_10_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_10_AWLEN <= twiddle_rsc_0_10_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_10_AWADDR <= twiddle_rsc_0_10_AWADDR;
  twiddle_rsc_0_11_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_11_RRESP;
  twiddle_rsc_0_11_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_11_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_11_ARREGION <= twiddle_rsc_0_11_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_11_ARQOS <= twiddle_rsc_0_11_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_11_ARPROT <= twiddle_rsc_0_11_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_11_ARCACHE <= twiddle_rsc_0_11_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_11_ARBURST <= twiddle_rsc_0_11_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_11_ARSIZE <= twiddle_rsc_0_11_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_11_ARLEN <= twiddle_rsc_0_11_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_11_ARADDR <= twiddle_rsc_0_11_ARADDR;
  twiddle_rsc_0_11_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_11_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_11_WSTRB <= twiddle_rsc_0_11_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_11_WDATA <= twiddle_rsc_0_11_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_11_AWREGION <= twiddle_rsc_0_11_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_11_AWQOS <= twiddle_rsc_0_11_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_11_AWPROT <= twiddle_rsc_0_11_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_11_AWCACHE <= twiddle_rsc_0_11_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_11_AWBURST <= twiddle_rsc_0_11_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_11_AWSIZE <= twiddle_rsc_0_11_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_11_AWLEN <= twiddle_rsc_0_11_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_11_AWADDR <= twiddle_rsc_0_11_AWADDR;
  twiddle_rsc_0_12_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_12_RRESP;
  twiddle_rsc_0_12_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_12_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_12_ARREGION <= twiddle_rsc_0_12_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_12_ARQOS <= twiddle_rsc_0_12_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_12_ARPROT <= twiddle_rsc_0_12_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_12_ARCACHE <= twiddle_rsc_0_12_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_12_ARBURST <= twiddle_rsc_0_12_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_12_ARSIZE <= twiddle_rsc_0_12_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_12_ARLEN <= twiddle_rsc_0_12_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_12_ARADDR <= twiddle_rsc_0_12_ARADDR;
  twiddle_rsc_0_12_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_12_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_12_WSTRB <= twiddle_rsc_0_12_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_12_WDATA <= twiddle_rsc_0_12_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_12_AWREGION <= twiddle_rsc_0_12_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_12_AWQOS <= twiddle_rsc_0_12_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_12_AWPROT <= twiddle_rsc_0_12_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_12_AWCACHE <= twiddle_rsc_0_12_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_12_AWBURST <= twiddle_rsc_0_12_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_12_AWSIZE <= twiddle_rsc_0_12_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_12_AWLEN <= twiddle_rsc_0_12_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_12_AWADDR <= twiddle_rsc_0_12_AWADDR;
  twiddle_rsc_0_13_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_13_RRESP;
  twiddle_rsc_0_13_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_13_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_13_ARREGION <= twiddle_rsc_0_13_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_13_ARQOS <= twiddle_rsc_0_13_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_13_ARPROT <= twiddle_rsc_0_13_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_13_ARCACHE <= twiddle_rsc_0_13_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_13_ARBURST <= twiddle_rsc_0_13_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_13_ARSIZE <= twiddle_rsc_0_13_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_13_ARLEN <= twiddle_rsc_0_13_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_13_ARADDR <= twiddle_rsc_0_13_ARADDR;
  twiddle_rsc_0_13_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_13_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_13_WSTRB <= twiddle_rsc_0_13_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_13_WDATA <= twiddle_rsc_0_13_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_13_AWREGION <= twiddle_rsc_0_13_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_13_AWQOS <= twiddle_rsc_0_13_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_13_AWPROT <= twiddle_rsc_0_13_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_13_AWCACHE <= twiddle_rsc_0_13_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_13_AWBURST <= twiddle_rsc_0_13_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_13_AWSIZE <= twiddle_rsc_0_13_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_13_AWLEN <= twiddle_rsc_0_13_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_13_AWADDR <= twiddle_rsc_0_13_AWADDR;
  twiddle_rsc_0_14_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_14_RRESP;
  twiddle_rsc_0_14_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_14_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_14_ARREGION <= twiddle_rsc_0_14_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_14_ARQOS <= twiddle_rsc_0_14_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_14_ARPROT <= twiddle_rsc_0_14_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_14_ARCACHE <= twiddle_rsc_0_14_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_14_ARBURST <= twiddle_rsc_0_14_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_14_ARSIZE <= twiddle_rsc_0_14_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_14_ARLEN <= twiddle_rsc_0_14_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_14_ARADDR <= twiddle_rsc_0_14_ARADDR;
  twiddle_rsc_0_14_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_14_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_14_WSTRB <= twiddle_rsc_0_14_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_14_WDATA <= twiddle_rsc_0_14_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_14_AWREGION <= twiddle_rsc_0_14_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_14_AWQOS <= twiddle_rsc_0_14_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_14_AWPROT <= twiddle_rsc_0_14_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_14_AWCACHE <= twiddle_rsc_0_14_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_14_AWBURST <= twiddle_rsc_0_14_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_14_AWSIZE <= twiddle_rsc_0_14_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_14_AWLEN <= twiddle_rsc_0_14_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_14_AWADDR <= twiddle_rsc_0_14_AWADDR;
  twiddle_rsc_0_15_RRESP <= peaseNTT_core_inst_twiddle_rsc_0_15_RRESP;
  twiddle_rsc_0_15_RDATA <= peaseNTT_core_inst_twiddle_rsc_0_15_RDATA;
  peaseNTT_core_inst_twiddle_rsc_0_15_ARREGION <= twiddle_rsc_0_15_ARREGION;
  peaseNTT_core_inst_twiddle_rsc_0_15_ARQOS <= twiddle_rsc_0_15_ARQOS;
  peaseNTT_core_inst_twiddle_rsc_0_15_ARPROT <= twiddle_rsc_0_15_ARPROT;
  peaseNTT_core_inst_twiddle_rsc_0_15_ARCACHE <= twiddle_rsc_0_15_ARCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_15_ARBURST <= twiddle_rsc_0_15_ARBURST;
  peaseNTT_core_inst_twiddle_rsc_0_15_ARSIZE <= twiddle_rsc_0_15_ARSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_15_ARLEN <= twiddle_rsc_0_15_ARLEN;
  peaseNTT_core_inst_twiddle_rsc_0_15_ARADDR <= twiddle_rsc_0_15_ARADDR;
  twiddle_rsc_0_15_BRESP <= peaseNTT_core_inst_twiddle_rsc_0_15_BRESP;
  peaseNTT_core_inst_twiddle_rsc_0_15_WSTRB <= twiddle_rsc_0_15_WSTRB;
  peaseNTT_core_inst_twiddle_rsc_0_15_WDATA <= twiddle_rsc_0_15_WDATA;
  peaseNTT_core_inst_twiddle_rsc_0_15_AWREGION <= twiddle_rsc_0_15_AWREGION;
  peaseNTT_core_inst_twiddle_rsc_0_15_AWQOS <= twiddle_rsc_0_15_AWQOS;
  peaseNTT_core_inst_twiddle_rsc_0_15_AWPROT <= twiddle_rsc_0_15_AWPROT;
  peaseNTT_core_inst_twiddle_rsc_0_15_AWCACHE <= twiddle_rsc_0_15_AWCACHE;
  peaseNTT_core_inst_twiddle_rsc_0_15_AWBURST <= twiddle_rsc_0_15_AWBURST;
  peaseNTT_core_inst_twiddle_rsc_0_15_AWSIZE <= twiddle_rsc_0_15_AWSIZE;
  peaseNTT_core_inst_twiddle_rsc_0_15_AWLEN <= twiddle_rsc_0_15_AWLEN;
  peaseNTT_core_inst_twiddle_rsc_0_15_AWADDR <= twiddle_rsc_0_15_AWADDR;
  twiddle_h_rsc_0_0_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_0_RRESP;
  twiddle_h_rsc_0_0_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_0_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_ARREGION <= twiddle_h_rsc_0_0_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_ARQOS <= twiddle_h_rsc_0_0_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_ARPROT <= twiddle_h_rsc_0_0_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_ARCACHE <= twiddle_h_rsc_0_0_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_ARBURST <= twiddle_h_rsc_0_0_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_ARSIZE <= twiddle_h_rsc_0_0_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_ARLEN <= twiddle_h_rsc_0_0_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_ARADDR <= twiddle_h_rsc_0_0_ARADDR;
  twiddle_h_rsc_0_0_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_0_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_WSTRB <= twiddle_h_rsc_0_0_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_WDATA <= twiddle_h_rsc_0_0_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_AWREGION <= twiddle_h_rsc_0_0_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_AWQOS <= twiddle_h_rsc_0_0_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_AWPROT <= twiddle_h_rsc_0_0_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_AWCACHE <= twiddle_h_rsc_0_0_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_AWBURST <= twiddle_h_rsc_0_0_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_AWSIZE <= twiddle_h_rsc_0_0_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_AWLEN <= twiddle_h_rsc_0_0_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_0_AWADDR <= twiddle_h_rsc_0_0_AWADDR;
  twiddle_h_rsc_0_1_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_1_RRESP;
  twiddle_h_rsc_0_1_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_1_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_ARREGION <= twiddle_h_rsc_0_1_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_ARQOS <= twiddle_h_rsc_0_1_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_ARPROT <= twiddle_h_rsc_0_1_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_ARCACHE <= twiddle_h_rsc_0_1_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_ARBURST <= twiddle_h_rsc_0_1_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_ARSIZE <= twiddle_h_rsc_0_1_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_ARLEN <= twiddle_h_rsc_0_1_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_ARADDR <= twiddle_h_rsc_0_1_ARADDR;
  twiddle_h_rsc_0_1_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_1_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_WSTRB <= twiddle_h_rsc_0_1_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_WDATA <= twiddle_h_rsc_0_1_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_AWREGION <= twiddle_h_rsc_0_1_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_AWQOS <= twiddle_h_rsc_0_1_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_AWPROT <= twiddle_h_rsc_0_1_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_AWCACHE <= twiddle_h_rsc_0_1_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_AWBURST <= twiddle_h_rsc_0_1_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_AWSIZE <= twiddle_h_rsc_0_1_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_AWLEN <= twiddle_h_rsc_0_1_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_1_AWADDR <= twiddle_h_rsc_0_1_AWADDR;
  twiddle_h_rsc_0_2_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_2_RRESP;
  twiddle_h_rsc_0_2_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_2_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_ARREGION <= twiddle_h_rsc_0_2_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_ARQOS <= twiddle_h_rsc_0_2_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_ARPROT <= twiddle_h_rsc_0_2_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_ARCACHE <= twiddle_h_rsc_0_2_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_ARBURST <= twiddle_h_rsc_0_2_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_ARSIZE <= twiddle_h_rsc_0_2_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_ARLEN <= twiddle_h_rsc_0_2_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_ARADDR <= twiddle_h_rsc_0_2_ARADDR;
  twiddle_h_rsc_0_2_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_2_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_WSTRB <= twiddle_h_rsc_0_2_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_WDATA <= twiddle_h_rsc_0_2_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_AWREGION <= twiddle_h_rsc_0_2_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_AWQOS <= twiddle_h_rsc_0_2_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_AWPROT <= twiddle_h_rsc_0_2_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_AWCACHE <= twiddle_h_rsc_0_2_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_AWBURST <= twiddle_h_rsc_0_2_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_AWSIZE <= twiddle_h_rsc_0_2_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_AWLEN <= twiddle_h_rsc_0_2_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_2_AWADDR <= twiddle_h_rsc_0_2_AWADDR;
  twiddle_h_rsc_0_3_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_3_RRESP;
  twiddle_h_rsc_0_3_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_3_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_ARREGION <= twiddle_h_rsc_0_3_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_ARQOS <= twiddle_h_rsc_0_3_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_ARPROT <= twiddle_h_rsc_0_3_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_ARCACHE <= twiddle_h_rsc_0_3_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_ARBURST <= twiddle_h_rsc_0_3_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_ARSIZE <= twiddle_h_rsc_0_3_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_ARLEN <= twiddle_h_rsc_0_3_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_ARADDR <= twiddle_h_rsc_0_3_ARADDR;
  twiddle_h_rsc_0_3_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_3_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_WSTRB <= twiddle_h_rsc_0_3_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_WDATA <= twiddle_h_rsc_0_3_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_AWREGION <= twiddle_h_rsc_0_3_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_AWQOS <= twiddle_h_rsc_0_3_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_AWPROT <= twiddle_h_rsc_0_3_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_AWCACHE <= twiddle_h_rsc_0_3_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_AWBURST <= twiddle_h_rsc_0_3_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_AWSIZE <= twiddle_h_rsc_0_3_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_AWLEN <= twiddle_h_rsc_0_3_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_3_AWADDR <= twiddle_h_rsc_0_3_AWADDR;
  twiddle_h_rsc_0_4_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_4_RRESP;
  twiddle_h_rsc_0_4_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_4_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_ARREGION <= twiddle_h_rsc_0_4_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_ARQOS <= twiddle_h_rsc_0_4_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_ARPROT <= twiddle_h_rsc_0_4_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_ARCACHE <= twiddle_h_rsc_0_4_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_ARBURST <= twiddle_h_rsc_0_4_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_ARSIZE <= twiddle_h_rsc_0_4_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_ARLEN <= twiddle_h_rsc_0_4_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_ARADDR <= twiddle_h_rsc_0_4_ARADDR;
  twiddle_h_rsc_0_4_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_4_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_WSTRB <= twiddle_h_rsc_0_4_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_WDATA <= twiddle_h_rsc_0_4_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_AWREGION <= twiddle_h_rsc_0_4_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_AWQOS <= twiddle_h_rsc_0_4_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_AWPROT <= twiddle_h_rsc_0_4_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_AWCACHE <= twiddle_h_rsc_0_4_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_AWBURST <= twiddle_h_rsc_0_4_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_AWSIZE <= twiddle_h_rsc_0_4_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_AWLEN <= twiddle_h_rsc_0_4_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_4_AWADDR <= twiddle_h_rsc_0_4_AWADDR;
  twiddle_h_rsc_0_5_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_5_RRESP;
  twiddle_h_rsc_0_5_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_5_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_ARREGION <= twiddle_h_rsc_0_5_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_ARQOS <= twiddle_h_rsc_0_5_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_ARPROT <= twiddle_h_rsc_0_5_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_ARCACHE <= twiddle_h_rsc_0_5_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_ARBURST <= twiddle_h_rsc_0_5_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_ARSIZE <= twiddle_h_rsc_0_5_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_ARLEN <= twiddle_h_rsc_0_5_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_ARADDR <= twiddle_h_rsc_0_5_ARADDR;
  twiddle_h_rsc_0_5_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_5_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_WSTRB <= twiddle_h_rsc_0_5_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_WDATA <= twiddle_h_rsc_0_5_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_AWREGION <= twiddle_h_rsc_0_5_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_AWQOS <= twiddle_h_rsc_0_5_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_AWPROT <= twiddle_h_rsc_0_5_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_AWCACHE <= twiddle_h_rsc_0_5_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_AWBURST <= twiddle_h_rsc_0_5_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_AWSIZE <= twiddle_h_rsc_0_5_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_AWLEN <= twiddle_h_rsc_0_5_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_5_AWADDR <= twiddle_h_rsc_0_5_AWADDR;
  twiddle_h_rsc_0_6_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_6_RRESP;
  twiddle_h_rsc_0_6_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_6_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_ARREGION <= twiddle_h_rsc_0_6_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_ARQOS <= twiddle_h_rsc_0_6_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_ARPROT <= twiddle_h_rsc_0_6_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_ARCACHE <= twiddle_h_rsc_0_6_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_ARBURST <= twiddle_h_rsc_0_6_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_ARSIZE <= twiddle_h_rsc_0_6_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_ARLEN <= twiddle_h_rsc_0_6_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_ARADDR <= twiddle_h_rsc_0_6_ARADDR;
  twiddle_h_rsc_0_6_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_6_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_WSTRB <= twiddle_h_rsc_0_6_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_WDATA <= twiddle_h_rsc_0_6_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_AWREGION <= twiddle_h_rsc_0_6_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_AWQOS <= twiddle_h_rsc_0_6_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_AWPROT <= twiddle_h_rsc_0_6_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_AWCACHE <= twiddle_h_rsc_0_6_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_AWBURST <= twiddle_h_rsc_0_6_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_AWSIZE <= twiddle_h_rsc_0_6_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_AWLEN <= twiddle_h_rsc_0_6_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_6_AWADDR <= twiddle_h_rsc_0_6_AWADDR;
  twiddle_h_rsc_0_7_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_7_RRESP;
  twiddle_h_rsc_0_7_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_7_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_ARREGION <= twiddle_h_rsc_0_7_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_ARQOS <= twiddle_h_rsc_0_7_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_ARPROT <= twiddle_h_rsc_0_7_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_ARCACHE <= twiddle_h_rsc_0_7_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_ARBURST <= twiddle_h_rsc_0_7_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_ARSIZE <= twiddle_h_rsc_0_7_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_ARLEN <= twiddle_h_rsc_0_7_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_ARADDR <= twiddle_h_rsc_0_7_ARADDR;
  twiddle_h_rsc_0_7_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_7_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_WSTRB <= twiddle_h_rsc_0_7_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_WDATA <= twiddle_h_rsc_0_7_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_AWREGION <= twiddle_h_rsc_0_7_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_AWQOS <= twiddle_h_rsc_0_7_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_AWPROT <= twiddle_h_rsc_0_7_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_AWCACHE <= twiddle_h_rsc_0_7_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_AWBURST <= twiddle_h_rsc_0_7_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_AWSIZE <= twiddle_h_rsc_0_7_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_AWLEN <= twiddle_h_rsc_0_7_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_7_AWADDR <= twiddle_h_rsc_0_7_AWADDR;
  twiddle_h_rsc_0_8_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_8_RRESP;
  twiddle_h_rsc_0_8_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_8_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_ARREGION <= twiddle_h_rsc_0_8_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_ARQOS <= twiddle_h_rsc_0_8_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_ARPROT <= twiddle_h_rsc_0_8_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_ARCACHE <= twiddle_h_rsc_0_8_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_ARBURST <= twiddle_h_rsc_0_8_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_ARSIZE <= twiddle_h_rsc_0_8_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_ARLEN <= twiddle_h_rsc_0_8_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_ARADDR <= twiddle_h_rsc_0_8_ARADDR;
  twiddle_h_rsc_0_8_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_8_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_WSTRB <= twiddle_h_rsc_0_8_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_WDATA <= twiddle_h_rsc_0_8_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_AWREGION <= twiddle_h_rsc_0_8_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_AWQOS <= twiddle_h_rsc_0_8_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_AWPROT <= twiddle_h_rsc_0_8_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_AWCACHE <= twiddle_h_rsc_0_8_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_AWBURST <= twiddle_h_rsc_0_8_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_AWSIZE <= twiddle_h_rsc_0_8_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_AWLEN <= twiddle_h_rsc_0_8_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_8_AWADDR <= twiddle_h_rsc_0_8_AWADDR;
  twiddle_h_rsc_0_9_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_9_RRESP;
  twiddle_h_rsc_0_9_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_9_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_ARREGION <= twiddle_h_rsc_0_9_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_ARQOS <= twiddle_h_rsc_0_9_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_ARPROT <= twiddle_h_rsc_0_9_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_ARCACHE <= twiddle_h_rsc_0_9_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_ARBURST <= twiddle_h_rsc_0_9_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_ARSIZE <= twiddle_h_rsc_0_9_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_ARLEN <= twiddle_h_rsc_0_9_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_ARADDR <= twiddle_h_rsc_0_9_ARADDR;
  twiddle_h_rsc_0_9_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_9_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_WSTRB <= twiddle_h_rsc_0_9_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_WDATA <= twiddle_h_rsc_0_9_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_AWREGION <= twiddle_h_rsc_0_9_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_AWQOS <= twiddle_h_rsc_0_9_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_AWPROT <= twiddle_h_rsc_0_9_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_AWCACHE <= twiddle_h_rsc_0_9_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_AWBURST <= twiddle_h_rsc_0_9_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_AWSIZE <= twiddle_h_rsc_0_9_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_AWLEN <= twiddle_h_rsc_0_9_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_9_AWADDR <= twiddle_h_rsc_0_9_AWADDR;
  twiddle_h_rsc_0_10_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_10_RRESP;
  twiddle_h_rsc_0_10_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_10_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_ARREGION <= twiddle_h_rsc_0_10_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_ARQOS <= twiddle_h_rsc_0_10_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_ARPROT <= twiddle_h_rsc_0_10_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_ARCACHE <= twiddle_h_rsc_0_10_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_ARBURST <= twiddle_h_rsc_0_10_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_ARSIZE <= twiddle_h_rsc_0_10_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_ARLEN <= twiddle_h_rsc_0_10_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_ARADDR <= twiddle_h_rsc_0_10_ARADDR;
  twiddle_h_rsc_0_10_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_10_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_WSTRB <= twiddle_h_rsc_0_10_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_WDATA <= twiddle_h_rsc_0_10_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_AWREGION <= twiddle_h_rsc_0_10_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_AWQOS <= twiddle_h_rsc_0_10_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_AWPROT <= twiddle_h_rsc_0_10_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_AWCACHE <= twiddle_h_rsc_0_10_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_AWBURST <= twiddle_h_rsc_0_10_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_AWSIZE <= twiddle_h_rsc_0_10_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_AWLEN <= twiddle_h_rsc_0_10_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_10_AWADDR <= twiddle_h_rsc_0_10_AWADDR;
  twiddle_h_rsc_0_11_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_11_RRESP;
  twiddle_h_rsc_0_11_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_11_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_ARREGION <= twiddle_h_rsc_0_11_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_ARQOS <= twiddle_h_rsc_0_11_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_ARPROT <= twiddle_h_rsc_0_11_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_ARCACHE <= twiddle_h_rsc_0_11_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_ARBURST <= twiddle_h_rsc_0_11_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_ARSIZE <= twiddle_h_rsc_0_11_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_ARLEN <= twiddle_h_rsc_0_11_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_ARADDR <= twiddle_h_rsc_0_11_ARADDR;
  twiddle_h_rsc_0_11_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_11_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_WSTRB <= twiddle_h_rsc_0_11_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_WDATA <= twiddle_h_rsc_0_11_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_AWREGION <= twiddle_h_rsc_0_11_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_AWQOS <= twiddle_h_rsc_0_11_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_AWPROT <= twiddle_h_rsc_0_11_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_AWCACHE <= twiddle_h_rsc_0_11_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_AWBURST <= twiddle_h_rsc_0_11_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_AWSIZE <= twiddle_h_rsc_0_11_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_AWLEN <= twiddle_h_rsc_0_11_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_11_AWADDR <= twiddle_h_rsc_0_11_AWADDR;
  twiddle_h_rsc_0_12_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_12_RRESP;
  twiddle_h_rsc_0_12_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_12_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_ARREGION <= twiddle_h_rsc_0_12_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_ARQOS <= twiddle_h_rsc_0_12_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_ARPROT <= twiddle_h_rsc_0_12_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_ARCACHE <= twiddle_h_rsc_0_12_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_ARBURST <= twiddle_h_rsc_0_12_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_ARSIZE <= twiddle_h_rsc_0_12_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_ARLEN <= twiddle_h_rsc_0_12_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_ARADDR <= twiddle_h_rsc_0_12_ARADDR;
  twiddle_h_rsc_0_12_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_12_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_WSTRB <= twiddle_h_rsc_0_12_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_WDATA <= twiddle_h_rsc_0_12_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_AWREGION <= twiddle_h_rsc_0_12_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_AWQOS <= twiddle_h_rsc_0_12_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_AWPROT <= twiddle_h_rsc_0_12_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_AWCACHE <= twiddle_h_rsc_0_12_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_AWBURST <= twiddle_h_rsc_0_12_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_AWSIZE <= twiddle_h_rsc_0_12_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_AWLEN <= twiddle_h_rsc_0_12_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_12_AWADDR <= twiddle_h_rsc_0_12_AWADDR;
  twiddle_h_rsc_0_13_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_13_RRESP;
  twiddle_h_rsc_0_13_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_13_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_ARREGION <= twiddle_h_rsc_0_13_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_ARQOS <= twiddle_h_rsc_0_13_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_ARPROT <= twiddle_h_rsc_0_13_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_ARCACHE <= twiddle_h_rsc_0_13_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_ARBURST <= twiddle_h_rsc_0_13_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_ARSIZE <= twiddle_h_rsc_0_13_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_ARLEN <= twiddle_h_rsc_0_13_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_ARADDR <= twiddle_h_rsc_0_13_ARADDR;
  twiddle_h_rsc_0_13_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_13_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_WSTRB <= twiddle_h_rsc_0_13_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_WDATA <= twiddle_h_rsc_0_13_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_AWREGION <= twiddle_h_rsc_0_13_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_AWQOS <= twiddle_h_rsc_0_13_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_AWPROT <= twiddle_h_rsc_0_13_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_AWCACHE <= twiddle_h_rsc_0_13_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_AWBURST <= twiddle_h_rsc_0_13_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_AWSIZE <= twiddle_h_rsc_0_13_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_AWLEN <= twiddle_h_rsc_0_13_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_13_AWADDR <= twiddle_h_rsc_0_13_AWADDR;
  twiddle_h_rsc_0_14_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_14_RRESP;
  twiddle_h_rsc_0_14_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_14_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_ARREGION <= twiddle_h_rsc_0_14_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_ARQOS <= twiddle_h_rsc_0_14_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_ARPROT <= twiddle_h_rsc_0_14_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_ARCACHE <= twiddle_h_rsc_0_14_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_ARBURST <= twiddle_h_rsc_0_14_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_ARSIZE <= twiddle_h_rsc_0_14_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_ARLEN <= twiddle_h_rsc_0_14_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_ARADDR <= twiddle_h_rsc_0_14_ARADDR;
  twiddle_h_rsc_0_14_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_14_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_WSTRB <= twiddle_h_rsc_0_14_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_WDATA <= twiddle_h_rsc_0_14_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_AWREGION <= twiddle_h_rsc_0_14_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_AWQOS <= twiddle_h_rsc_0_14_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_AWPROT <= twiddle_h_rsc_0_14_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_AWCACHE <= twiddle_h_rsc_0_14_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_AWBURST <= twiddle_h_rsc_0_14_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_AWSIZE <= twiddle_h_rsc_0_14_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_AWLEN <= twiddle_h_rsc_0_14_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_14_AWADDR <= twiddle_h_rsc_0_14_AWADDR;
  twiddle_h_rsc_0_15_RRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_15_RRESP;
  twiddle_h_rsc_0_15_RDATA <= peaseNTT_core_inst_twiddle_h_rsc_0_15_RDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_ARREGION <= twiddle_h_rsc_0_15_ARREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_ARQOS <= twiddle_h_rsc_0_15_ARQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_ARPROT <= twiddle_h_rsc_0_15_ARPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_ARCACHE <= twiddle_h_rsc_0_15_ARCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_ARBURST <= twiddle_h_rsc_0_15_ARBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_ARSIZE <= twiddle_h_rsc_0_15_ARSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_ARLEN <= twiddle_h_rsc_0_15_ARLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_ARADDR <= twiddle_h_rsc_0_15_ARADDR;
  twiddle_h_rsc_0_15_BRESP <= peaseNTT_core_inst_twiddle_h_rsc_0_15_BRESP;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_WSTRB <= twiddle_h_rsc_0_15_WSTRB;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_WDATA <= twiddle_h_rsc_0_15_WDATA;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_AWREGION <= twiddle_h_rsc_0_15_AWREGION;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_AWQOS <= twiddle_h_rsc_0_15_AWQOS;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_AWPROT <= twiddle_h_rsc_0_15_AWPROT;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_AWCACHE <= twiddle_h_rsc_0_15_AWCACHE;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_AWBURST <= twiddle_h_rsc_0_15_AWBURST;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_AWSIZE <= twiddle_h_rsc_0_15_AWSIZE;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_AWLEN <= twiddle_h_rsc_0_15_AWLEN;
  peaseNTT_core_inst_twiddle_h_rsc_0_15_AWADDR <= twiddle_h_rsc_0_15_AWADDR;
  peaseNTT_core_inst_yt_rsc_0_0_i_qa_d <= yt_rsc_0_0_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_1_i_qa_d <= yt_rsc_0_1_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_2_i_qa_d <= yt_rsc_0_2_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_3_i_qa_d <= yt_rsc_0_3_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_4_i_qa_d <= yt_rsc_0_4_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_5_i_qa_d <= yt_rsc_0_5_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_6_i_qa_d <= yt_rsc_0_6_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_7_i_qa_d <= yt_rsc_0_7_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_8_i_qa_d <= yt_rsc_0_8_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_9_i_qa_d <= yt_rsc_0_9_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_10_i_qa_d <= yt_rsc_0_10_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_11_i_qa_d <= yt_rsc_0_11_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_12_i_qa_d <= yt_rsc_0_12_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_13_i_qa_d <= yt_rsc_0_13_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_14_i_qa_d <= yt_rsc_0_14_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_15_i_qa_d <= yt_rsc_0_15_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_16_i_qa_d <= yt_rsc_0_16_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_17_i_qa_d <= yt_rsc_0_17_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_18_i_qa_d <= yt_rsc_0_18_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_19_i_qa_d <= yt_rsc_0_19_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_20_i_qa_d <= yt_rsc_0_20_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_21_i_qa_d <= yt_rsc_0_21_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_22_i_qa_d <= yt_rsc_0_22_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_23_i_qa_d <= yt_rsc_0_23_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_24_i_qa_d <= yt_rsc_0_24_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_25_i_qa_d <= yt_rsc_0_25_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_26_i_qa_d <= yt_rsc_0_26_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_27_i_qa_d <= yt_rsc_0_27_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_28_i_qa_d <= yt_rsc_0_28_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_29_i_qa_d <= yt_rsc_0_29_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_30_i_qa_d <= yt_rsc_0_30_i_qa_d;
  peaseNTT_core_inst_yt_rsc_0_31_i_qa_d <= yt_rsc_0_31_i_qa_d;
  yt_rsc_1_0_i_da_d <= peaseNTT_core_inst_yt_rsc_1_0_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_0_i_qa_d <= yt_rsc_1_0_i_qa_d;
  yt_rsc_1_1_i_da_d <= peaseNTT_core_inst_yt_rsc_1_1_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_1_i_qa_d <= yt_rsc_1_1_i_qa_d;
  yt_rsc_1_2_i_da_d <= peaseNTT_core_inst_yt_rsc_1_2_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_2_i_qa_d <= yt_rsc_1_2_i_qa_d;
  yt_rsc_1_3_i_da_d <= peaseNTT_core_inst_yt_rsc_1_3_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_3_i_qa_d <= yt_rsc_1_3_i_qa_d;
  yt_rsc_1_4_i_da_d <= peaseNTT_core_inst_yt_rsc_1_4_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_4_i_qa_d <= yt_rsc_1_4_i_qa_d;
  yt_rsc_1_5_i_da_d <= peaseNTT_core_inst_yt_rsc_1_5_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_5_i_qa_d <= yt_rsc_1_5_i_qa_d;
  yt_rsc_1_6_i_da_d <= peaseNTT_core_inst_yt_rsc_1_6_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_6_i_qa_d <= yt_rsc_1_6_i_qa_d;
  yt_rsc_1_7_i_da_d <= peaseNTT_core_inst_yt_rsc_1_7_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_7_i_qa_d <= yt_rsc_1_7_i_qa_d;
  yt_rsc_1_8_i_da_d <= peaseNTT_core_inst_yt_rsc_1_8_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_8_i_qa_d <= yt_rsc_1_8_i_qa_d;
  yt_rsc_1_9_i_da_d <= peaseNTT_core_inst_yt_rsc_1_9_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_9_i_qa_d <= yt_rsc_1_9_i_qa_d;
  yt_rsc_1_10_i_da_d <= peaseNTT_core_inst_yt_rsc_1_10_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_10_i_qa_d <= yt_rsc_1_10_i_qa_d;
  yt_rsc_1_11_i_da_d <= peaseNTT_core_inst_yt_rsc_1_11_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_11_i_qa_d <= yt_rsc_1_11_i_qa_d;
  yt_rsc_1_12_i_da_d <= peaseNTT_core_inst_yt_rsc_1_12_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_12_i_qa_d <= yt_rsc_1_12_i_qa_d;
  yt_rsc_1_13_i_da_d <= peaseNTT_core_inst_yt_rsc_1_13_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_13_i_qa_d <= yt_rsc_1_13_i_qa_d;
  yt_rsc_1_14_i_da_d <= peaseNTT_core_inst_yt_rsc_1_14_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_14_i_qa_d <= yt_rsc_1_14_i_qa_d;
  yt_rsc_1_15_i_da_d <= peaseNTT_core_inst_yt_rsc_1_15_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_15_i_qa_d <= yt_rsc_1_15_i_qa_d;
  yt_rsc_1_16_i_da_d <= peaseNTT_core_inst_yt_rsc_1_16_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_16_i_qa_d <= yt_rsc_1_16_i_qa_d;
  yt_rsc_1_17_i_da_d <= peaseNTT_core_inst_yt_rsc_1_17_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_17_i_qa_d <= yt_rsc_1_17_i_qa_d;
  yt_rsc_1_18_i_da_d <= peaseNTT_core_inst_yt_rsc_1_18_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_18_i_qa_d <= yt_rsc_1_18_i_qa_d;
  yt_rsc_1_19_i_da_d <= peaseNTT_core_inst_yt_rsc_1_19_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_19_i_qa_d <= yt_rsc_1_19_i_qa_d;
  yt_rsc_1_20_i_da_d <= peaseNTT_core_inst_yt_rsc_1_20_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_20_i_qa_d <= yt_rsc_1_20_i_qa_d;
  yt_rsc_1_21_i_da_d <= peaseNTT_core_inst_yt_rsc_1_21_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_21_i_qa_d <= yt_rsc_1_21_i_qa_d;
  yt_rsc_1_22_i_da_d <= peaseNTT_core_inst_yt_rsc_1_22_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_22_i_qa_d <= yt_rsc_1_22_i_qa_d;
  yt_rsc_1_23_i_da_d <= peaseNTT_core_inst_yt_rsc_1_23_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_23_i_qa_d <= yt_rsc_1_23_i_qa_d;
  yt_rsc_1_24_i_da_d <= peaseNTT_core_inst_yt_rsc_1_24_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_24_i_qa_d <= yt_rsc_1_24_i_qa_d;
  yt_rsc_1_25_i_da_d <= peaseNTT_core_inst_yt_rsc_1_25_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_25_i_qa_d <= yt_rsc_1_25_i_qa_d;
  yt_rsc_1_26_i_da_d <= peaseNTT_core_inst_yt_rsc_1_26_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_26_i_qa_d <= yt_rsc_1_26_i_qa_d;
  yt_rsc_1_27_i_da_d <= peaseNTT_core_inst_yt_rsc_1_27_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_27_i_qa_d <= yt_rsc_1_27_i_qa_d;
  yt_rsc_1_28_i_da_d <= peaseNTT_core_inst_yt_rsc_1_28_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_28_i_qa_d <= yt_rsc_1_28_i_qa_d;
  yt_rsc_1_29_i_da_d <= peaseNTT_core_inst_yt_rsc_1_29_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_29_i_qa_d <= yt_rsc_1_29_i_qa_d;
  yt_rsc_1_30_i_da_d <= peaseNTT_core_inst_yt_rsc_1_30_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_30_i_qa_d <= yt_rsc_1_30_i_qa_d;
  yt_rsc_1_31_i_da_d <= peaseNTT_core_inst_yt_rsc_1_31_i_da_d;
  peaseNTT_core_inst_yt_rsc_1_31_i_qa_d <= yt_rsc_1_31_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_0_i_qa_d <= xt_rsc_0_0_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_1_i_qa_d <= xt_rsc_0_1_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_2_i_qa_d <= xt_rsc_0_2_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_3_i_qa_d <= xt_rsc_0_3_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_4_i_qa_d <= xt_rsc_0_4_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_5_i_qa_d <= xt_rsc_0_5_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_6_i_qa_d <= xt_rsc_0_6_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_7_i_qa_d <= xt_rsc_0_7_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_8_i_qa_d <= xt_rsc_0_8_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_9_i_qa_d <= xt_rsc_0_9_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_10_i_qa_d <= xt_rsc_0_10_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_11_i_qa_d <= xt_rsc_0_11_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_12_i_qa_d <= xt_rsc_0_12_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_13_i_qa_d <= xt_rsc_0_13_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_14_i_qa_d <= xt_rsc_0_14_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_15_i_qa_d <= xt_rsc_0_15_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_16_i_qa_d <= xt_rsc_0_16_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_17_i_qa_d <= xt_rsc_0_17_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_18_i_qa_d <= xt_rsc_0_18_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_19_i_qa_d <= xt_rsc_0_19_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_20_i_qa_d <= xt_rsc_0_20_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_21_i_qa_d <= xt_rsc_0_21_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_22_i_qa_d <= xt_rsc_0_22_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_23_i_qa_d <= xt_rsc_0_23_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_24_i_qa_d <= xt_rsc_0_24_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_25_i_qa_d <= xt_rsc_0_25_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_26_i_qa_d <= xt_rsc_0_26_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_27_i_qa_d <= xt_rsc_0_27_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_28_i_qa_d <= xt_rsc_0_28_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_29_i_qa_d <= xt_rsc_0_29_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_30_i_qa_d <= xt_rsc_0_30_i_qa_d;
  peaseNTT_core_inst_xt_rsc_0_31_i_qa_d <= xt_rsc_0_31_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_0_i_qa_d <= xt_rsc_1_0_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_1_i_qa_d <= xt_rsc_1_1_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_2_i_qa_d <= xt_rsc_1_2_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_3_i_qa_d <= xt_rsc_1_3_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_4_i_qa_d <= xt_rsc_1_4_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_5_i_qa_d <= xt_rsc_1_5_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_6_i_qa_d <= xt_rsc_1_6_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_7_i_qa_d <= xt_rsc_1_7_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_8_i_qa_d <= xt_rsc_1_8_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_9_i_qa_d <= xt_rsc_1_9_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_10_i_qa_d <= xt_rsc_1_10_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_11_i_qa_d <= xt_rsc_1_11_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_12_i_qa_d <= xt_rsc_1_12_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_13_i_qa_d <= xt_rsc_1_13_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_14_i_qa_d <= xt_rsc_1_14_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_15_i_qa_d <= xt_rsc_1_15_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_16_i_qa_d <= xt_rsc_1_16_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_17_i_qa_d <= xt_rsc_1_17_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_18_i_qa_d <= xt_rsc_1_18_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_19_i_qa_d <= xt_rsc_1_19_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_20_i_qa_d <= xt_rsc_1_20_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_21_i_qa_d <= xt_rsc_1_21_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_22_i_qa_d <= xt_rsc_1_22_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_23_i_qa_d <= xt_rsc_1_23_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_24_i_qa_d <= xt_rsc_1_24_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_25_i_qa_d <= xt_rsc_1_25_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_26_i_qa_d <= xt_rsc_1_26_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_27_i_qa_d <= xt_rsc_1_27_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_28_i_qa_d <= xt_rsc_1_28_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_29_i_qa_d <= xt_rsc_1_29_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_30_i_qa_d <= xt_rsc_1_30_i_qa_d;
  peaseNTT_core_inst_xt_rsc_1_31_i_qa_d <= xt_rsc_1_31_i_qa_d;
  yt_rsc_0_0_i_adra_d_iff <= peaseNTT_core_inst_yt_rsc_0_0_i_adra_d_pff;
  yt_rsc_0_0_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_0_i_da_d_pff;
  yt_rsc_0_1_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_1_i_da_d_pff;
  yt_rsc_0_2_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_2_i_da_d_pff;
  yt_rsc_0_3_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_3_i_da_d_pff;
  yt_rsc_0_4_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_4_i_da_d_pff;
  yt_rsc_0_5_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_5_i_da_d_pff;
  yt_rsc_0_6_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_6_i_da_d_pff;
  yt_rsc_0_7_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_7_i_da_d_pff;
  yt_rsc_0_8_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_8_i_da_d_pff;
  yt_rsc_0_9_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_9_i_da_d_pff;
  yt_rsc_0_10_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_10_i_da_d_pff;
  yt_rsc_0_11_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_11_i_da_d_pff;
  yt_rsc_0_12_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_12_i_da_d_pff;
  yt_rsc_0_13_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_13_i_da_d_pff;
  yt_rsc_0_14_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_14_i_da_d_pff;
  yt_rsc_0_15_i_da_d_iff <= peaseNTT_core_inst_yt_rsc_0_15_i_da_d_pff;
  yt_rsc_0_16_i_adra_d_iff <= peaseNTT_core_inst_yt_rsc_0_16_i_adra_d_pff;
  yt_rsc_1_0_i_adra_d_iff <= peaseNTT_core_inst_yt_rsc_1_0_i_adra_d_pff;
  yt_rsc_1_16_i_adra_d_iff <= peaseNTT_core_inst_yt_rsc_1_16_i_adra_d_pff;
  xt_rsc_0_0_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_0_i_adra_d_pff;
  xt_rsc_0_0_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_0_i_da_d_pff;
  xt_rsc_0_1_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_1_i_da_d_pff;
  xt_rsc_0_2_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_2_i_da_d_pff;
  xt_rsc_0_3_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_3_i_da_d_pff;
  xt_rsc_0_4_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_4_i_da_d_pff;
  xt_rsc_0_5_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_5_i_da_d_pff;
  xt_rsc_0_6_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_6_i_da_d_pff;
  xt_rsc_0_7_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_7_i_da_d_pff;
  xt_rsc_0_8_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_8_i_da_d_pff;
  xt_rsc_0_9_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_9_i_da_d_pff;
  xt_rsc_0_10_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_10_i_da_d_pff;
  xt_rsc_0_11_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_11_i_da_d_pff;
  xt_rsc_0_12_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_12_i_da_d_pff;
  xt_rsc_0_13_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_13_i_da_d_pff;
  xt_rsc_0_14_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_14_i_da_d_pff;
  xt_rsc_0_15_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_0_15_i_da_d_pff;
  xt_rsc_0_16_i_adra_d_iff <= peaseNTT_core_inst_xt_rsc_0_16_i_adra_d_pff;
  xt_rsc_1_0_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_0_i_da_d_pff;
  xt_rsc_1_1_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_1_i_da_d_pff;
  xt_rsc_1_2_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_2_i_da_d_pff;
  xt_rsc_1_3_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_3_i_da_d_pff;
  xt_rsc_1_4_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_4_i_da_d_pff;
  xt_rsc_1_5_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_5_i_da_d_pff;
  xt_rsc_1_6_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_6_i_da_d_pff;
  xt_rsc_1_7_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_7_i_da_d_pff;
  xt_rsc_1_8_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_8_i_da_d_pff;
  xt_rsc_1_9_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_9_i_da_d_pff;
  xt_rsc_1_10_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_10_i_da_d_pff;
  xt_rsc_1_11_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_11_i_da_d_pff;
  xt_rsc_1_12_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_12_i_da_d_pff;
  xt_rsc_1_13_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_13_i_da_d_pff;
  xt_rsc_1_14_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_14_i_da_d_pff;
  xt_rsc_1_15_i_da_d_iff <= peaseNTT_core_inst_xt_rsc_1_15_i_da_d_pff;

END v29;



