
//------> /opt/mentorgraphics/Catapult_10.3a/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/mentorgraphics/Catapult_10.3a/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /opt/mentorgraphics/Catapult_10.3a/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.3a/798110 Production Release
//  HLS Date:       Tue Dec  4 22:20:19 PST 2018
// 
//  Generated by:   jd4691@newnano.poly.edu
//  Generated date: Wed Jun 23 00:11:20 2021
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_filter_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module fir_filter_core_core_fsm (
  clk, rst, fsm_output, SHIFT_LOOP_C_0_tr0, MAC_LOOP_C_0_tr0
);
  input clk;
  input rst;
  output [4:0] fsm_output;
  reg [4:0] fsm_output;
  input SHIFT_LOOP_C_0_tr0;
  input MAC_LOOP_C_0_tr0;


  // FSM State Type Declaration for fir_filter_core_core_fsm_1
  parameter
    main_C_0 = 3'd0,
    SHIFT_LOOP_C_0 = 3'd1,
    MAC_LOOP_C_0 = 3'd2,
    main_C_1 = 3'd3,
    main_C_2 = 3'd4;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : fir_filter_core_core_fsm_1
    case (state_var)
      SHIFT_LOOP_C_0 : begin
        fsm_output = 5'b00010;
        if ( SHIFT_LOOP_C_0_tr0 ) begin
          state_var_NS = MAC_LOOP_C_0;
        end
        else begin
          state_var_NS = SHIFT_LOOP_C_0;
        end
      end
      MAC_LOOP_C_0 : begin
        fsm_output = 5'b00100;
        if ( MAC_LOOP_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = MAC_LOOP_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 5'b01000;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 5'b10000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 5'b00001;
        state_var_NS = SHIFT_LOOP_C_0;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_filter_core
// ------------------------------------------------------------------


module fir_filter_core (
  clk, rst, i_sample_rsc_dat, i_sample_rsc_triosy_lz, b_rsc_dat, b_rsc_triosy_lz,
      y_rsc_dat, y_rsc_triosy_lz
);
  input clk;
  input rst;
  input [2:0] i_sample_rsc_dat;
  output i_sample_rsc_triosy_lz;
  input [1269:0] b_rsc_dat;
  output b_rsc_triosy_lz;
  output [8:0] y_rsc_dat;
  output y_rsc_triosy_lz;


  // Interconnect Declarations
  wire [2:0] i_sample_rsci_idat;
  wire [1269:0] b_rsci_idat;
  reg y_rsc_triosy_obj_ld;
  reg y_rsci_idat_8;
  reg [6:0] y_rsci_idat_7_1;
  reg y_rsci_idat_0;
  wire [4:0] fsm_output;
  reg [6:0] MAC_LOOP_n_6_0_sva;
  reg [19:0] sum_sva;
  reg reg_b_rsc_triosy_obj_ld_cse;
  wire [2:0] z_out;
  wire [19:0] z_out_2;
  wire [20:0] nl_z_out_2;
  reg [2:0] x_0_sva;
  reg [2:0] x_63_lpi_2;
  reg [2:0] x_62_lpi_2;
  reg [2:0] x_64_lpi_2;
  reg [2:0] x_61_lpi_2;
  reg [2:0] x_65_lpi_2;
  reg [2:0] x_60_lpi_2;
  reg [2:0] x_66_lpi_2;
  reg [2:0] x_59_lpi_2;
  reg [2:0] x_67_lpi_2;
  reg [2:0] x_58_lpi_2;
  reg [2:0] x_68_lpi_2;
  reg [2:0] x_57_lpi_2;
  reg [2:0] x_69_lpi_2;
  reg [2:0] x_56_lpi_2;
  reg [2:0] x_70_lpi_2;
  reg [2:0] x_55_lpi_2;
  reg [2:0] x_71_lpi_2;
  reg [2:0] x_54_lpi_2;
  reg [2:0] x_72_lpi_2;
  reg [2:0] x_53_lpi_2;
  reg [2:0] x_73_lpi_2;
  reg [2:0] x_52_lpi_2;
  reg [2:0] x_74_lpi_2;
  reg [2:0] x_51_lpi_2;
  reg [2:0] x_75_lpi_2;
  reg [2:0] x_50_lpi_2;
  reg [2:0] x_76_lpi_2;
  reg [2:0] x_49_lpi_2;
  reg [2:0] x_77_lpi_2;
  reg [2:0] x_48_lpi_2;
  reg [2:0] x_78_lpi_2;
  reg [2:0] x_47_lpi_2;
  reg [2:0] x_79_lpi_2;
  reg [2:0] x_46_lpi_2;
  reg [2:0] x_80_lpi_2;
  reg [2:0] x_45_lpi_2;
  reg [2:0] x_81_lpi_2;
  reg [2:0] x_44_lpi_2;
  reg [2:0] x_82_lpi_2;
  reg [2:0] x_43_lpi_2;
  reg [2:0] x_83_lpi_2;
  reg [2:0] x_42_lpi_2;
  reg [2:0] x_84_lpi_2;
  reg [2:0] x_41_lpi_2;
  reg [2:0] x_85_lpi_2;
  reg [2:0] x_40_lpi_2;
  reg [2:0] x_86_lpi_2;
  reg [2:0] x_39_lpi_2;
  reg [2:0] x_87_lpi_2;
  reg [2:0] x_38_lpi_2;
  reg [2:0] x_88_lpi_2;
  reg [2:0] x_37_lpi_2;
  reg [2:0] x_89_lpi_2;
  reg [2:0] x_36_lpi_2;
  reg [2:0] x_90_lpi_2;
  reg [2:0] x_35_lpi_2;
  reg [2:0] x_91_lpi_2;
  reg [2:0] x_34_lpi_2;
  reg [2:0] x_92_lpi_2;
  reg [2:0] x_33_lpi_2;
  reg [2:0] x_93_lpi_2;
  reg [2:0] x_32_lpi_2;
  reg [2:0] x_94_lpi_2;
  reg [2:0] x_31_lpi_2;
  reg [2:0] x_95_lpi_2;
  reg [2:0] x_30_lpi_2;
  reg [2:0] x_96_lpi_2;
  reg [2:0] x_29_lpi_2;
  reg [2:0] x_97_lpi_2;
  reg [2:0] x_28_lpi_2;
  reg [2:0] x_98_lpi_2;
  reg [2:0] x_27_lpi_2;
  reg [2:0] x_99_lpi_2;
  reg [2:0] x_26_lpi_2;
  reg [2:0] x_100_lpi_2;
  reg [2:0] x_25_lpi_2;
  reg [2:0] x_101_lpi_2;
  reg [2:0] x_24_lpi_2;
  reg [2:0] x_102_lpi_2;
  reg [2:0] x_23_lpi_2;
  reg [2:0] x_103_lpi_2;
  reg [2:0] x_22_lpi_2;
  reg [2:0] x_104_lpi_2;
  reg [2:0] x_21_lpi_2;
  reg [2:0] x_105_lpi_2;
  reg [2:0] x_20_lpi_2;
  reg [2:0] x_106_lpi_2;
  reg [2:0] x_19_lpi_2;
  reg [2:0] x_107_lpi_2;
  reg [2:0] x_18_lpi_2;
  reg [2:0] x_108_lpi_2;
  reg [2:0] x_17_lpi_2;
  reg [2:0] x_109_lpi_2;
  reg [2:0] x_16_lpi_2;
  reg [2:0] x_110_lpi_2;
  reg [2:0] x_15_lpi_2;
  reg [2:0] x_111_lpi_2;
  reg [2:0] x_14_lpi_2;
  reg [2:0] x_112_lpi_2;
  reg [2:0] x_13_lpi_2;
  reg [2:0] x_113_lpi_2;
  reg [2:0] x_12_lpi_2;
  reg [2:0] x_114_lpi_2;
  reg [2:0] x_11_lpi_2;
  reg [2:0] x_115_lpi_2;
  reg [2:0] x_10_lpi_2;
  reg [2:0] x_116_lpi_2;
  reg [2:0] x_9_lpi_2;
  reg [2:0] x_117_lpi_2;
  reg [2:0] x_8_lpi_2;
  reg [2:0] x_118_lpi_2;
  reg [2:0] x_7_lpi_2;
  reg [2:0] x_119_lpi_2;
  reg [2:0] x_6_lpi_2;
  reg [2:0] x_120_lpi_2;
  reg [2:0] x_5_lpi_2;
  reg [2:0] x_121_lpi_2;
  reg [2:0] x_4_lpi_2;
  reg [2:0] x_122_lpi_2;
  reg [2:0] x_3_lpi_2;
  reg [2:0] x_123_lpi_2;
  reg [2:0] x_2_lpi_2;
  reg [2:0] x_124_lpi_2;
  reg [2:0] x_1_lpi_2;
  reg [2:0] x_125_lpi_2;
  reg [2:0] x_126_lpi_2;
  reg [2:0] i_sample_sva;
  wire nor_ovfl_sva_1;
  wire and_unfl_sva_1;
  wire z_out_1_7;
  wire [6:0] MAC_LOOP_mux_11_tmp;
  wire and_tmp;
  wire and_tmp_2;
  wire and_tmp_3;
  wire and_tmp_5;
  wire and_tmp_6;
  wire and_tmp_7;
  wire and_tmp_8;
  wire and_tmp_9;
  wire and_tmp_10;
  wire and_tmp_12;
  wire and_tmp_13;
  wire and_tmp_14;
  wire and_tmp_15;
  wire and_tmp_16;
  wire and_tmp_17;
  wire and_tmp_18;
  wire and_tmp_19;
  wire and_tmp_20;
  wire and_tmp_21;
  wire and_tmp_22;
  wire and_tmp_23;
  wire and_tmp_24;
  wire and_tmp_25;
  wire and_tmp_26;
  wire and_tmp_27;
  wire and_tmp_28;
  wire and_tmp_29;
  wire and_tmp_30;
  wire and_tmp_31;
  wire and_tmp_32;
  wire and_tmp_33;
  wire and_tmp_34;
  wire and_tmp_35;
  wire and_tmp_36;
  wire and_tmp_37;
  wire and_tmp_38;
  wire and_tmp_39;
  wire and_tmp_40;
  wire and_tmp_41;
  wire and_tmp_42;
  wire and_tmp_43;
  wire and_tmp_44;
  wire and_tmp_45;
  wire and_tmp_46;
  wire and_tmp_47;
  wire and_tmp_48;
  wire and_tmp_49;
  wire and_tmp_50;
  wire and_tmp_51;
  wire and_tmp_52;
  wire and_tmp_53;
  wire and_tmp_54;
  wire and_tmp_55;
  wire and_tmp_56;
  wire and_tmp_57;
  wire and_tmp_58;
  wire and_tmp_59;
  wire and_tmp_60;
  wire and_tmp_61;
  wire and_tmp_62;
  wire and_tmp_63;
  wire and_tmp_64;
  wire and_tmp_65;
  wire and_tmp_66;
  wire and_tmp_67;
  wire and_tmp_68;
  wire and_tmp_69;
  wire and_tmp_70;
  wire and_tmp_71;
  wire and_tmp_72;
  wire and_tmp_73;
  wire and_tmp_74;
  wire and_tmp_75;
  wire and_tmp_76;
  wire and_tmp_77;
  wire and_tmp_78;
  wire and_tmp_79;
  wire and_tmp_80;
  wire and_tmp_81;
  wire and_tmp_82;
  wire and_tmp_83;
  wire and_tmp_84;
  wire and_tmp_85;
  wire and_tmp_86;
  wire and_tmp_87;
  wire and_tmp_88;
  wire and_tmp_89;
  wire and_tmp_90;
  wire and_tmp_91;
  wire and_tmp_92;
  wire and_tmp_93;
  wire and_tmp_94;
  wire and_tmp_95;
  wire and_tmp_96;
  wire and_tmp_97;
  wire and_tmp_98;
  wire and_tmp_99;
  wire and_tmp_100;
  wire and_tmp_101;
  wire and_tmp_102;
  wire and_tmp_103;
  wire and_tmp_104;
  wire and_tmp_105;
  wire and_tmp_106;
  wire and_tmp_107;
  wire and_tmp_108;
  wire and_tmp_109;
  wire and_tmp_110;
  wire and_tmp_111;
  wire and_tmp_112;
  wire and_tmp_113;
  wire and_tmp_114;
  wire and_tmp_115;
  wire and_tmp_116;
  wire and_tmp_117;
  wire and_tmp_118;
  wire [6:0] acc_2_tmp_7_1;
  wire [7:0] nl_acc_2_tmp_7_1;
  wire nor_1308_cse;
  wire nor_1309_cse;
  wire and_2671_cse;
  wire and_2667_cse;
  wire nor_1303_cse;
  wire and_2691_cse;
  wire and_2736_cse;
  wire and_2741_cse;
  wire and_2829_cse;
  wire nor_1310_cse;
  wire and_2668_cse;
  wire nor_1297_cse;
  wire and_2677_cse;
  wire nor_1259_cse;
  wire and_2708_cse;
  wire nor_1271_cse;
  wire and_2698_cse;
  wire nor_1240_cse;
  wire and_2723_cse;
  wire nor_1202_cse;
  wire and_2753_cse;
  wire nor_1184_cse;
  wire and_2768_cse;
  wire nor_1188_cse;
  wire and_2765_cse;
  wire nor_1213_cse;
  wire and_2743_cse;
  wire nor_1159_cse;
  wire and_2792_cse;
  wire nor_1149_cse;
  wire and_2801_cse;
  wire nor_1132_cse;
  wire and_2816_cse;
  wire nor_1098_cse;
  wire and_2846_cse;
  wire nor_1077_cse;
  wire and_2861_cse;
  wire nor_1082_cse;
  wire and_2858_cse;
  wire nor_1048_cse;
  wire and_2885_cse;
  wire nor_1037_cse;
  wire and_2894_cse;
  wire nor_1052_cse;
  wire and_2882_cse;
  wire nor_1017_cse;
  wire and_2909_cse;
  wire nor_986_cse;
  wire and_2933_cse;
  wire nor_975_cse;
  wire and_2942_cse;
  wire nor_956_cse;
  wire and_2957_cse;
  wire nor_960_cse;
  wire and_2954_cse;
  wire nor_931_cse;
  wire and_2981_cse;
  wire nor_921_cse;
  wire and_2990_cse;
  wire nor_905_cse;
  wire and_3005_cse;

  wire[6:0] nor_5_nl;
  wire[0:0] mux_221_nl;
  wire[0:0] nor_1306_nl;
  wire[0:0] nor_1307_nl;
  wire[0:0] mux_222_nl;
  wire[0:0] mux_224_nl;
  wire[0:0] nor_1299_nl;
  wire[0:0] nor_1300_nl;
  wire[0:0] mux_226_nl;
  wire[0:0] nor_1293_nl;
  wire[0:0] nor_1294_nl;
  wire[0:0] mux_227_nl;
  wire[0:0] mux_229_nl;
  wire[0:0] nor_1287_nl;
  wire[0:0] nor_1288_nl;
  wire[0:0] mux_231_nl;
  wire[0:0] nor_1285_nl;
  wire[0:0] nor_1286_nl;
  wire[0:0] mux_233_nl;
  wire[0:0] nor_1281_nl;
  wire[0:0] nor_1282_nl;
  wire[0:0] mux_235_nl;
  wire[0:0] nor_1278_nl;
  wire[0:0] nor_1279_nl;
  wire[0:0] mux_237_nl;
  wire[0:0] nor_1273_nl;
  wire[0:0] nor_1274_nl;
  wire[0:0] mux_239_nl;
  wire[0:0] nor_1268_nl;
  wire[0:0] nor_1269_nl;
  wire[0:0] mux_240_nl;
  wire[0:0] mux_242_nl;
  wire[0:0] nor_1262_nl;
  wire[0:0] nor_1263_nl;
  wire[0:0] mux_244_nl;
  wire[0:0] nor_1260_nl;
  wire[0:0] nor_1261_nl;
  wire[0:0] mux_246_nl;
  wire[0:0] nor_1256_nl;
  wire[0:0] nor_1257_nl;
  wire[0:0] mux_248_nl;
  wire[0:0] nor_1253_nl;
  wire[0:0] nor_1254_nl;
  wire[0:0] mux_250_nl;
  wire[0:0] nor_1248_nl;
  wire[0:0] nor_1249_nl;
  wire[0:0] mux_252_nl;
  wire[0:0] nor_1245_nl;
  wire[0:0] nor_1246_nl;
  wire[0:0] mux_254_nl;
  wire[0:0] nor_1241_nl;
  wire[0:0] nor_1242_nl;
  wire[0:0] mux_256_nl;
  wire[0:0] nor_1237_nl;
  wire[0:0] nor_1238_nl;
  wire[0:0] mux_258_nl;
  wire[0:0] nor_1232_nl;
  wire[0:0] nor_1233_nl;
  wire[0:0] mux_260_nl;
  wire[0:0] nor_1228_nl;
  wire[0:0] nor_1229_nl;
  wire[0:0] mux_262_nl;
  wire[0:0] nor_1224_nl;
  wire[0:0] nor_1225_nl;
  wire[0:0] mux_264_nl;
  wire[0:0] nor_1220_nl;
  wire[0:0] nor_1221_nl;
  wire[0:0] mux_266_nl;
  wire[0:0] nor_1215_nl;
  wire[0:0] nor_1216_nl;
  wire[0:0] mux_268_nl;
  wire[0:0] nor_1210_nl;
  wire[0:0] nor_1211_nl;
  wire[0:0] mux_270_nl;
  wire[0:0] or_1206_nl;
  wire[0:0] mux_272_nl;
  wire[0:0] nor_1205_nl;
  wire[0:0] nor_1206_nl;
  wire[0:0] mux_274_nl;
  wire[0:0] nor_1203_nl;
  wire[0:0] nor_1204_nl;
  wire[0:0] mux_276_nl;
  wire[0:0] nor_1199_nl;
  wire[0:0] nor_1200_nl;
  wire[0:0] mux_278_nl;
  wire[0:0] nor_1196_nl;
  wire[0:0] nor_1197_nl;
  wire[0:0] mux_280_nl;
  wire[0:0] nor_1191_nl;
  wire[0:0] nor_1192_nl;
  wire[0:0] mux_282_nl;
  wire[0:0] nor_1189_nl;
  wire[0:0] nor_1190_nl;
  wire[0:0] mux_284_nl;
  wire[0:0] nor_1185_nl;
  wire[0:0] nor_1186_nl;
  wire[0:0] mux_286_nl;
  wire[0:0] nor_1182_nl;
  wire[0:0] nor_1183_nl;
  wire[0:0] mux_288_nl;
  wire[0:0] nor_1178_nl;
  wire[0:0] nor_1179_nl;
  wire[0:0] mux_290_nl;
  wire[0:0] nor_1175_nl;
  wire[0:0] nor_1176_nl;
  wire[0:0] mux_292_nl;
  wire[0:0] nor_1172_nl;
  wire[0:0] nor_1173_nl;
  wire[0:0] mux_294_nl;
  wire[0:0] nor_1169_nl;
  wire[0:0] nor_1170_nl;
  wire[0:0] mux_296_nl;
  wire[0:0] nor_1165_nl;
  wire[0:0] nor_1166_nl;
  wire[0:0] mux_298_nl;
  wire[0:0] nor_1163_nl;
  wire[0:0] nor_1164_nl;
  wire[0:0] mux_300_nl;
  wire[0:0] nor_1160_nl;
  wire[0:0] nor_1161_nl;
  wire[0:0] mux_302_nl;
  wire[0:0] nor_1157_nl;
  wire[0:0] nor_1158_nl;
  wire[0:0] mux_304_nl;
  wire[0:0] nor_1153_nl;
  wire[0:0] nor_1154_nl;
  wire[0:0] mux_306_nl;
  wire[0:0] nor_1150_nl;
  wire[0:0] nor_1151_nl;
  wire[0:0] mux_308_nl;
  wire[0:0] nor_1147_nl;
  wire[0:0] nor_1148_nl;
  wire[0:0] mux_310_nl;
  wire[0:0] nor_1144_nl;
  wire[0:0] nor_1145_nl;
  wire[0:0] mux_312_nl;
  wire[0:0] nor_1140_nl;
  wire[0:0] nor_1141_nl;
  wire[0:0] mux_314_nl;
  wire[0:0] nor_1136_nl;
  wire[0:0] nor_1137_nl;
  wire[0:0] mux_316_nl;
  wire[0:0] nor_1133_nl;
  wire[0:0] nor_1134_nl;
  wire[0:0] mux_318_nl;
  wire[0:0] nor_1129_nl;
  wire[0:0] nor_1130_nl;
  wire[0:0] mux_320_nl;
  wire[0:0] nor_1125_nl;
  wire[0:0] nor_1126_nl;
  wire[0:0] mux_322_nl;
  wire[0:0] nor_1121_nl;
  wire[0:0] nor_1122_nl;
  wire[0:0] mux_324_nl;
  wire[0:0] nor_1118_nl;
  wire[0:0] nor_1119_nl;
  wire[0:0] mux_326_nl;
  wire[0:0] nor_1114_nl;
  wire[0:0] nor_1115_nl;
  wire[0:0] mux_328_nl;
  wire[0:0] nor_1110_nl;
  wire[0:0] nor_1111_nl;
  wire[0:0] mux_330_nl;
  wire[0:0] nor_1107_nl;
  wire[0:0] nor_1108_nl;
  wire[0:0] mux_332_nl;
  wire[0:0] or_1205_nl;
  wire[0:0] mux_334_nl;
  wire[0:0] nor_1101_nl;
  wire[0:0] nor_1102_nl;
  wire[0:0] mux_336_nl;
  wire[0:0] nor_1099_nl;
  wire[0:0] nor_1100_nl;
  wire[0:0] mux_338_nl;
  wire[0:0] nor_1094_nl;
  wire[0:0] nor_1095_nl;
  wire[0:0] mux_340_nl;
  wire[0:0] nor_1090_nl;
  wire[0:0] nor_1091_nl;
  wire[0:0] mux_342_nl;
  wire[0:0] nor_1085_nl;
  wire[0:0] nor_1086_nl;
  wire[0:0] mux_344_nl;
  wire[0:0] nor_1083_nl;
  wire[0:0] nor_1084_nl;
  wire[0:0] mux_346_nl;
  wire[0:0] nor_1078_nl;
  wire[0:0] nor_1079_nl;
  wire[0:0] mux_348_nl;
  wire[0:0] nor_1074_nl;
  wire[0:0] nor_1075_nl;
  wire[0:0] mux_350_nl;
  wire[0:0] nor_1070_nl;
  wire[0:0] nor_1071_nl;
  wire[0:0] mux_352_nl;
  wire[0:0] nor_1067_nl;
  wire[0:0] nor_1068_nl;
  wire[0:0] mux_354_nl;
  wire[0:0] nor_1063_nl;
  wire[0:0] nor_1064_nl;
  wire[0:0] mux_356_nl;
  wire[0:0] nor_1059_nl;
  wire[0:0] nor_1060_nl;
  wire[0:0] mux_358_nl;
  wire[0:0] nor_1055_nl;
  wire[0:0] nor_1056_nl;
  wire[0:0] mux_360_nl;
  wire[0:0] nor_1053_nl;
  wire[0:0] nor_1054_nl;
  wire[0:0] mux_362_nl;
  wire[0:0] nor_1049_nl;
  wire[0:0] nor_1050_nl;
  wire[0:0] mux_364_nl;
  wire[0:0] nor_1045_nl;
  wire[0:0] nor_1046_nl;
  wire[0:0] mux_366_nl;
  wire[0:0] nor_1041_nl;
  wire[0:0] nor_1042_nl;
  wire[0:0] mux_368_nl;
  wire[0:0] nor_1038_nl;
  wire[0:0] nor_1039_nl;
  wire[0:0] mux_370_nl;
  wire[0:0] nor_1034_nl;
  wire[0:0] nor_1035_nl;
  wire[0:0] mux_372_nl;
  wire[0:0] nor_1030_nl;
  wire[0:0] nor_1031_nl;
  wire[0:0] mux_374_nl;
  wire[0:0] nor_1026_nl;
  wire[0:0] nor_1027_nl;
  wire[0:0] mux_376_nl;
  wire[0:0] nor_1022_nl;
  wire[0:0] nor_1023_nl;
  wire[0:0] mux_378_nl;
  wire[0:0] nor_1018_nl;
  wire[0:0] nor_1019_nl;
  wire[0:0] mux_380_nl;
  wire[0:0] nor_1013_nl;
  wire[0:0] nor_1014_nl;
  wire[0:0] mux_382_nl;
  wire[0:0] nor_1009_nl;
  wire[0:0] nor_1010_nl;
  wire[0:0] mux_384_nl;
  wire[0:0] nor_1005_nl;
  wire[0:0] nor_1006_nl;
  wire[0:0] mux_386_nl;
  wire[0:0] nor_1001_nl;
  wire[0:0] nor_1002_nl;
  wire[0:0] mux_388_nl;
  wire[0:0] nor_996_nl;
  wire[0:0] nor_997_nl;
  wire[0:0] mux_390_nl;
  wire[0:0] nor_992_nl;
  wire[0:0] nor_993_nl;
  wire[0:0] mux_392_nl;
  wire[0:0] nor_990_nl;
  wire[0:0] nor_991_nl;
  wire[0:0] mux_394_nl;
  wire[0:0] nor_987_nl;
  wire[0:0] nor_988_nl;
  wire[0:0] mux_396_nl;
  wire[0:0] nor_983_nl;
  wire[0:0] nor_984_nl;
  wire[0:0] mux_398_nl;
  wire[0:0] nor_979_nl;
  wire[0:0] nor_980_nl;
  wire[0:0] mux_400_nl;
  wire[0:0] nor_976_nl;
  wire[0:0] nor_977_nl;
  wire[0:0] mux_402_nl;
  wire[0:0] nor_972_nl;
  wire[0:0] nor_973_nl;
  wire[0:0] mux_404_nl;
  wire[0:0] nor_968_nl;
  wire[0:0] nor_969_nl;
  wire[0:0] mux_406_nl;
  wire[0:0] nor_964_nl;
  wire[0:0] nor_965_nl;
  wire[0:0] mux_408_nl;
  wire[0:0] nor_961_nl;
  wire[0:0] nor_962_nl;
  wire[0:0] mux_410_nl;
  wire[0:0] nor_957_nl;
  wire[0:0] nor_958_nl;
  wire[0:0] mux_412_nl;
  wire[0:0] nor_953_nl;
  wire[0:0] nor_954_nl;
  wire[0:0] mux_414_nl;
  wire[0:0] nor_950_nl;
  wire[0:0] nor_951_nl;
  wire[0:0] mux_416_nl;
  wire[0:0] nor_947_nl;
  wire[0:0] nor_948_nl;
  wire[0:0] mux_418_nl;
  wire[0:0] nor_944_nl;
  wire[0:0] nor_945_nl;
  wire[0:0] mux_420_nl;
  wire[0:0] nor_940_nl;
  wire[0:0] nor_941_nl;
  wire[0:0] mux_422_nl;
  wire[0:0] nor_937_nl;
  wire[0:0] nor_938_nl;
  wire[0:0] mux_424_nl;
  wire[0:0] nor_934_nl;
  wire[0:0] nor_935_nl;
  wire[0:0] mux_426_nl;
  wire[0:0] nor_932_nl;
  wire[0:0] nor_933_nl;
  wire[0:0] mux_428_nl;
  wire[0:0] nor_928_nl;
  wire[0:0] nor_929_nl;
  wire[0:0] mux_430_nl;
  wire[0:0] nor_925_nl;
  wire[0:0] nor_926_nl;
  wire[0:0] mux_432_nl;
  wire[0:0] nor_922_nl;
  wire[0:0] nor_923_nl;
  wire[0:0] mux_434_nl;
  wire[0:0] nor_919_nl;
  wire[0:0] nor_920_nl;
  wire[0:0] mux_436_nl;
  wire[0:0] nor_915_nl;
  wire[0:0] nor_916_nl;
  wire[0:0] mux_438_nl;
  wire[0:0] nor_912_nl;
  wire[0:0] nor_913_nl;
  wire[0:0] mux_440_nl;
  wire[0:0] nor_908_nl;
  wire[0:0] nor_909_nl;
  wire[0:0] mux_442_nl;
  wire[0:0] nor_906_nl;
  wire[0:0] nor_907_nl;
  wire[0:0] mux_444_nl;
  wire[0:0] nor_901_nl;
  wire[0:0] nor_902_nl;
  wire[0:0] mux_446_nl;
  wire[0:0] nor_898_nl;
  wire[0:0] nor_899_nl;
  wire[0:0] mux_448_nl;
  wire[0:0] nor_894_nl;
  wire[0:0] nor_895_nl;
  wire[0:0] mux_450_nl;
  wire[0:0] nor_892_nl;
  wire[0:0] nor_893_nl;
  wire[0:0] mux_452_nl;
  wire[0:0] nor_887_nl;
  wire[0:0] nor_888_nl;
  wire[0:0] mux_454_nl;
  wire[0:0] or_1204_nl;
  wire[6:0] SHIFT_LOOP_n_SHIFT_LOOP_n_mux_nl;
  wire[0:0] SHIFT_LOOP_n_or_nl;
  wire[0:0] MAC_LOOP_n_nor_nl;
  wire[0:0] mux_220_nl;
  wire[0:0] mux_223_nl;
  wire[0:0] mux_225_nl;
  wire[0:0] mux_228_nl;
  wire[0:0] nor_1291_nl;
  wire[0:0] and_2681_nl;
  wire[0:0] mux_230_nl;
  wire[0:0] mux_232_nl;
  wire[0:0] mux_234_nl;
  wire[0:0] nor_1280_nl;
  wire[0:0] and_2690_nl;
  wire[0:0] mux_236_nl;
  wire[0:0] mux_238_nl;
  wire[0:0] mux_241_nl;
  wire[0:0] nor_1266_nl;
  wire[0:0] and_2702_nl;
  wire[0:0] mux_243_nl;
  wire[0:0] mux_245_nl;
  wire[0:0] mux_247_nl;
  wire[0:0] nor_1255_nl;
  wire[0:0] and_2711_nl;
  wire[0:0] mux_249_nl;
  wire[0:0] mux_251_nl;
  wire[0:0] mux_253_nl;
  wire[0:0] mux_255_nl;
  wire[0:0] mux_257_nl;
  wire[0:0] nor_1236_nl;
  wire[0:0] and_2726_nl;
  wire[0:0] mux_259_nl;
  wire[0:0] mux_261_nl;
  wire[0:0] mux_263_nl;
  wire[0:0] nor_1223_nl;
  wire[0:0] and_2735_nl;
  wire[0:0] mux_265_nl;
  wire[0:0] mux_267_nl;
  wire[0:0] mux_269_nl;
  wire[0:0] mux_271_nl;
  wire[0:0] nor_1209_nl;
  wire[0:0] and_2747_nl;
  wire[0:0] mux_273_nl;
  wire[0:0] mux_275_nl;
  wire[0:0] mux_277_nl;
  wire[0:0] nor_1198_nl;
  wire[0:0] and_2756_nl;
  wire[0:0] mux_279_nl;
  wire[0:0] mux_281_nl;
  wire[0:0] mux_283_nl;
  wire[0:0] mux_285_nl;
  wire[0:0] mux_287_nl;
  wire[0:0] nor_1181_nl;
  wire[0:0] and_2771_nl;
  wire[0:0] mux_289_nl;
  wire[0:0] mux_291_nl;
  wire[0:0] mux_293_nl;
  wire[0:0] nor_1171_nl;
  wire[0:0] and_2780_nl;
  wire[0:0] mux_295_nl;
  wire[0:0] mux_297_nl;
  wire[0:0] mux_299_nl;
  wire[0:0] mux_301_nl;
  wire[0:0] mux_303_nl;
  wire[0:0] nor_1156_nl;
  wire[0:0] and_2795_nl;
  wire[0:0] mux_305_nl;
  wire[0:0] mux_307_nl;
  wire[0:0] mux_309_nl;
  wire[0:0] nor_1146_nl;
  wire[0:0] and_2804_nl;
  wire[0:0] mux_311_nl;
  wire[0:0] mux_313_nl;
  wire[0:0] mux_315_nl;
  wire[0:0] mux_317_nl;
  wire[0:0] mux_319_nl;
  wire[0:0] nor_1128_nl;
  wire[0:0] and_2819_nl;
  wire[0:0] mux_321_nl;
  wire[0:0] mux_323_nl;
  wire[0:0] mux_325_nl;
  wire[0:0] nor_1117_nl;
  wire[0:0] and_2828_nl;
  wire[0:0] mux_327_nl;
  wire[0:0] mux_329_nl;
  wire[0:0] mux_331_nl;
  wire[0:0] mux_333_nl;
  wire[0:0] nor_1105_nl;
  wire[0:0] and_2840_nl;
  wire[0:0] mux_335_nl;
  wire[0:0] mux_337_nl;
  wire[0:0] mux_339_nl;
  wire[0:0] nor_1093_nl;
  wire[0:0] and_2849_nl;
  wire[0:0] mux_341_nl;
  wire[0:0] mux_343_nl;
  wire[0:0] mux_345_nl;
  wire[0:0] mux_347_nl;
  wire[0:0] mux_349_nl;
  wire[0:0] nor_1073_nl;
  wire[0:0] and_2864_nl;
  wire[0:0] mux_351_nl;
  wire[0:0] mux_353_nl;
  wire[0:0] mux_355_nl;
  wire[0:0] nor_1062_nl;
  wire[0:0] and_2873_nl;
  wire[0:0] mux_357_nl;
  wire[0:0] mux_359_nl;
  wire[0:0] mux_361_nl;
  wire[0:0] mux_363_nl;
  wire[0:0] mux_365_nl;
  wire[0:0] nor_1044_nl;
  wire[0:0] and_2888_nl;
  wire[0:0] mux_367_nl;
  wire[0:0] mux_369_nl;
  wire[0:0] mux_371_nl;
  wire[0:0] nor_1033_nl;
  wire[0:0] and_2897_nl;
  wire[0:0] mux_373_nl;
  wire[0:0] mux_375_nl;
  wire[0:0] mux_377_nl;
  wire[0:0] mux_379_nl;
  wire[0:0] mux_381_nl;
  wire[0:0] nor_1012_nl;
  wire[0:0] and_2912_nl;
  wire[0:0] mux_383_nl;
  wire[0:0] mux_385_nl;
  wire[0:0] mux_387_nl;
  wire[0:0] nor_1000_nl;
  wire[0:0] and_2921_nl;
  wire[0:0] mux_389_nl;
  wire[0:0] mux_391_nl;
  wire[0:0] mux_393_nl;
  wire[0:0] mux_395_nl;
  wire[0:0] mux_397_nl;
  wire[0:0] nor_982_nl;
  wire[0:0] and_2936_nl;
  wire[0:0] mux_399_nl;
  wire[0:0] mux_401_nl;
  wire[0:0] mux_403_nl;
  wire[0:0] nor_971_nl;
  wire[0:0] and_2945_nl;
  wire[0:0] mux_405_nl;
  wire[0:0] mux_407_nl;
  wire[0:0] mux_409_nl;
  wire[0:0] mux_411_nl;
  wire[0:0] mux_413_nl;
  wire[0:0] nor_952_nl;
  wire[0:0] and_2960_nl;
  wire[0:0] mux_415_nl;
  wire[0:0] mux_417_nl;
  wire[0:0] mux_419_nl;
  wire[0:0] nor_943_nl;
  wire[0:0] and_2969_nl;
  wire[0:0] mux_421_nl;
  wire[0:0] mux_423_nl;
  wire[0:0] mux_425_nl;
  wire[0:0] mux_427_nl;
  wire[0:0] mux_429_nl;
  wire[0:0] nor_927_nl;
  wire[0:0] and_2984_nl;
  wire[0:0] mux_431_nl;
  wire[0:0] mux_433_nl;
  wire[0:0] mux_435_nl;
  wire[0:0] nor_918_nl;
  wire[0:0] and_2993_nl;
  wire[0:0] mux_437_nl;
  wire[0:0] mux_439_nl;
  wire[0:0] mux_441_nl;
  wire[0:0] mux_443_nl;
  wire[0:0] mux_445_nl;
  wire[0:0] nor_900_nl;
  wire[0:0] and_3008_nl;
  wire[0:0] mux_447_nl;
  wire[0:0] mux_449_nl;
  wire[0:0] mux_451_nl;
  wire[0:0] nor_891_nl;
  wire[0:0] and_3016_nl;
  wire[0:0] mux_453_nl;
  wire[7:0] SHIFT_LOOP_acc_nl;
  wire[8:0] nl_SHIFT_LOOP_acc_nl;
  wire[6:0] SHIFT_LOOP_mux_129_nl;
  wire[18:0] MAC_LOOP_mux_7_nl;
  wire[12:0] MAC_LOOP_mux_8_nl;
  wire[12:0] MAC_LOOP_mul_1_nl;
  wire[9:0] MAC_LOOP_mux_9_nl;
  wire[2:0] MAC_LOOP_mux_10_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [8:0] nl_y_rsci_idat;
  assign nl_y_rsci_idat = {y_rsci_idat_8 , y_rsci_idat_7_1 , y_rsci_idat_0};
  wire [0:0] nl_fir_filter_core_core_fsm_inst_SHIFT_LOOP_C_0_tr0;
  assign nl_fir_filter_core_core_fsm_inst_SHIFT_LOOP_C_0_tr0 = ~ z_out_1_7;
  wire [0:0] nl_fir_filter_core_core_fsm_inst_MAC_LOOP_C_0_tr0;
  assign nl_fir_filter_core_core_fsm_inst_MAC_LOOP_C_0_tr0 = ~ z_out_1_7;
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd3)) i_sample_rsci (
      .dat(i_sample_rsc_dat),
      .idat(i_sample_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd1270)) b_rsci (
      .dat(b_rsc_dat),
      .idat(b_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd3),
  .width(32'sd9)) y_rsci (
      .idat(nl_y_rsci_idat[8:0]),
      .dat(y_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) i_sample_rsc_triosy_obj (
      .ld(reg_b_rsc_triosy_obj_ld_cse),
      .lz(i_sample_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) b_rsc_triosy_obj (
      .ld(reg_b_rsc_triosy_obj_ld_cse),
      .lz(b_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) y_rsc_triosy_obj (
      .ld(y_rsc_triosy_obj_ld),
      .lz(y_rsc_triosy_lz)
    );
  fir_filter_core_core_fsm fir_filter_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output),
      .SHIFT_LOOP_C_0_tr0(nl_fir_filter_core_core_fsm_inst_SHIFT_LOOP_C_0_tr0[0:0]),
      .MAC_LOOP_C_0_tr0(nl_fir_filter_core_core_fsm_inst_MAC_LOOP_C_0_tr0[0:0])
    );
  assign nor_1308_cse = ~((MAC_LOOP_n_6_0_sva[3:2]!=2'b00));
  assign nor_1309_cse = ~((MAC_LOOP_n_6_0_sva[4]) | (MAC_LOOP_n_6_0_sva[6]));
  assign and_2667_cse = (acc_2_tmp_7_1[6:2]==5'b11111);
  assign and_2671_cse = (acc_2_tmp_7_1[3]) & (acc_2_tmp_7_1[4]) & (acc_2_tmp_7_1[5])
      & (acc_2_tmp_7_1[6]) & (acc_2_tmp_7_1[1]);
  assign nor_1303_cse = ~((MAC_LOOP_n_6_0_sva[5]) | (MAC_LOOP_n_6_0_sva[0]));
  assign and_2691_cse = (acc_2_tmp_7_1[4]) & (acc_2_tmp_7_1[5]) & (acc_2_tmp_7_1[6])
      & (acc_2_tmp_7_1[1]) & (acc_2_tmp_7_1[2]);
  assign and_2736_cse = (acc_2_tmp_7_1[5]) & (acc_2_tmp_7_1[6]) & (acc_2_tmp_7_1[3])
      & (acc_2_tmp_7_1[2]) & (acc_2_tmp_7_1[1]);
  assign and_2741_cse = (acc_2_tmp_7_1[5:1]==5'b11111);
  assign and_2829_cse = (acc_2_tmp_7_1[6]) & (acc_2_tmp_7_1[4]) & (acc_2_tmp_7_1[3])
      & (acc_2_tmp_7_1[2]) & (acc_2_tmp_7_1[1]);
  assign nor_ovfl_sva_1 = ~((z_out_2[14]) | (~((z_out_2[13:8]!=6'b000000))));
  assign and_unfl_sva_1 = (z_out_2[14]) & (~((z_out_2[13:8]==6'b111111) & ((z_out_2[7:0]!=8'b00000000))));
  assign nor_1310_cse = ~((MAC_LOOP_mux_11_tmp[6:2]!=5'b00000));
  assign and_2668_cse = (MAC_LOOP_mux_11_tmp[6:2]==5'b11111);
  assign mux_220_nl = MUX_s_1_2_2(nor_1310_cse, and_2668_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp = (MAC_LOOP_mux_11_tmp[0]) & (mux_220_nl);
  assign mux_223_nl = MUX_s_1_2_2(nor_1310_cse, and_2668_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_2 = (MAC_LOOP_mux_11_tmp[1]) & (mux_223_nl);
  assign nor_1297_cse = ~((MAC_LOOP_mux_11_tmp[6:3]!=4'b0000));
  assign and_2677_cse = (MAC_LOOP_mux_11_tmp[6:3]==4'b1111);
  assign mux_225_nl = MUX_s_1_2_2(nor_1297_cse, and_2677_cse, MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_3 = (MAC_LOOP_mux_11_tmp[1:0]==2'b11) & (mux_225_nl);
  assign nor_1291_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[4])
      | (MAC_LOOP_mux_11_tmp[5]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2681_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_228_nl = MUX_s_1_2_2((nor_1291_nl), (and_2681_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_5 = (MAC_LOOP_mux_11_tmp[2]) & (mux_228_nl);
  assign mux_230_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[2])), (MAC_LOOP_mux_11_tmp[2]),
      MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_6 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_230_nl);
  assign mux_232_nl = MUX_s_1_2_2(nor_1297_cse, and_2677_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_7 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (mux_232_nl);
  assign nor_1280_nl = ~((MAC_LOOP_mux_11_tmp[2:1]!=2'b00));
  assign and_2690_nl = (MAC_LOOP_mux_11_tmp[2:1]==2'b11);
  assign mux_234_nl = MUX_s_1_2_2((nor_1280_nl), (and_2690_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_8 = (MAC_LOOP_mux_11_tmp[6:3]==4'b1111) & (mux_234_nl);
  assign mux_236_nl = MUX_s_1_2_2(nor_1297_cse, and_2677_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_9 = (MAC_LOOP_mux_11_tmp[2:1]==2'b11) & (mux_236_nl);
  assign nor_1271_cse = ~((MAC_LOOP_mux_11_tmp[6:4]!=3'b000));
  assign and_2698_cse = (MAC_LOOP_mux_11_tmp[6:4]==3'b111);
  assign mux_238_nl = MUX_s_1_2_2(nor_1271_cse, and_2698_cse, MAC_LOOP_mux_11_tmp[3]);
  assign and_tmp_10 = (MAC_LOOP_mux_11_tmp[2:0]==3'b111) & (mux_238_nl);
  assign nor_1266_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[4])
      | (MAC_LOOP_mux_11_tmp[5]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2702_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_241_nl = MUX_s_1_2_2((nor_1266_nl), (and_2702_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_12 = (MAC_LOOP_mux_11_tmp[3]) & (mux_241_nl);
  assign mux_243_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[3])), (MAC_LOOP_mux_11_tmp[3]),
      MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_13 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_243_nl);
  assign nor_1259_cse = ~((MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[4]) | (MAC_LOOP_mux_11_tmp[5])
      | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2708_cse = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5])
      & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_245_nl = MUX_s_1_2_2(nor_1259_cse, and_2708_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_14 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[3]) & (mux_245_nl);
  assign nor_1255_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[3]));
  assign and_2711_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]);
  assign mux_247_nl = MUX_s_1_2_2((nor_1255_nl), (and_2711_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_15 = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_247_nl);
  assign mux_249_nl = MUX_s_1_2_2(nor_1259_cse, and_2708_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_16 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (mux_249_nl);
  assign mux_251_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[3])), (MAC_LOOP_mux_11_tmp[3]),
      MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_17 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_251_nl);
  assign mux_253_nl = MUX_s_1_2_2(nor_1271_cse, and_2698_cse, MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_18 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3])
      & (mux_253_nl);
  assign nor_1240_cse = ~((MAC_LOOP_mux_11_tmp[3:2]!=2'b00));
  assign and_2723_cse = (MAC_LOOP_mux_11_tmp[3:2]==2'b11);
  assign mux_255_nl = MUX_s_1_2_2(nor_1240_cse, and_2723_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_19 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_255_nl);
  assign nor_1236_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[4]) | (MAC_LOOP_mux_11_tmp[5])
      | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2726_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5])
      & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_257_nl = MUX_s_1_2_2((nor_1236_nl), (and_2726_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_20 = (MAC_LOOP_mux_11_tmp[3:2]==2'b11) & (mux_257_nl);
  assign mux_259_nl = MUX_s_1_2_2(nor_1240_cse, and_2723_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_21 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_259_nl);
  assign mux_261_nl = MUX_s_1_2_2(nor_1271_cse, and_2698_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_22 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (mux_261_nl);
  assign nor_1223_nl = ~((MAC_LOOP_mux_11_tmp[3:1]!=3'b000));
  assign and_2735_nl = (MAC_LOOP_mux_11_tmp[3:1]==3'b111);
  assign mux_263_nl = MUX_s_1_2_2((nor_1223_nl), (and_2735_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_23 = (MAC_LOOP_mux_11_tmp[6:4]==3'b111) & (mux_263_nl);
  assign mux_265_nl = MUX_s_1_2_2(nor_1271_cse, and_2698_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_24 = (MAC_LOOP_mux_11_tmp[3:1]==3'b111) & (mux_265_nl);
  assign nor_1213_cse = ~((MAC_LOOP_mux_11_tmp[6:5]!=2'b00));
  assign and_2743_cse = (MAC_LOOP_mux_11_tmp[6:5]==2'b11);
  assign mux_267_nl = MUX_s_1_2_2(nor_1213_cse, and_2743_cse, MAC_LOOP_mux_11_tmp[4]);
  assign and_tmp_25 = (MAC_LOOP_mux_11_tmp[3:0]==4'b1111) & (mux_267_nl);
  assign mux_269_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[4])), (MAC_LOOP_mux_11_tmp[4]),
      MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_26 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_269_nl);
  assign nor_1209_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[3])
      | (MAC_LOOP_mux_11_tmp[5]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2747_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_271_nl = MUX_s_1_2_2((nor_1209_nl), (and_2747_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_27 = (MAC_LOOP_mux_11_tmp[4]) & (mux_271_nl);
  assign mux_273_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[4])), (MAC_LOOP_mux_11_tmp[4]),
      MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_28 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_273_nl);
  assign nor_1202_cse = ~((MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[5])
      | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2753_cse = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5])
      & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_275_nl = MUX_s_1_2_2(nor_1202_cse, and_2753_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_29 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[4]) & (mux_275_nl);
  assign nor_1198_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[4]));
  assign and_2756_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[4]);
  assign mux_277_nl = MUX_s_1_2_2((nor_1198_nl), (and_2756_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_30 = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_277_nl);
  assign mux_279_nl = MUX_s_1_2_2(nor_1202_cse, and_2753_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_31 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[4]) & (mux_279_nl);
  assign mux_281_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[4])), (MAC_LOOP_mux_11_tmp[4]),
      MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_32 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_281_nl);
  assign nor_1188_cse = ~((MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[5]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2765_cse = (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_283_nl = MUX_s_1_2_2(nor_1188_cse, and_2765_cse, MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_33 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[4])
      & (mux_283_nl);
  assign nor_1184_cse = ~((MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[4]));
  assign and_2768_cse = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4]);
  assign mux_285_nl = MUX_s_1_2_2(nor_1184_cse, and_2768_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_34 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_285_nl);
  assign nor_1181_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[5])
      | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2771_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5])
      & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_287_nl = MUX_s_1_2_2((nor_1181_nl), (and_2771_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_35 = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4]) & (mux_287_nl);
  assign mux_289_nl = MUX_s_1_2_2(nor_1184_cse, and_2768_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_36 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_289_nl);
  assign mux_291_nl = MUX_s_1_2_2(nor_1188_cse, and_2765_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_37 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4])
      & (mux_291_nl);
  assign nor_1171_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[4]));
  assign and_2780_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4]);
  assign mux_293_nl = MUX_s_1_2_2((nor_1171_nl), (and_2780_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_38 = (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6])
      & (mux_293_nl);
  assign mux_295_nl = MUX_s_1_2_2(nor_1188_cse, and_2765_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_39 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4])
      & (mux_295_nl);
  assign mux_297_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[4])), (MAC_LOOP_mux_11_tmp[4]),
      MAC_LOOP_mux_11_tmp[3]);
  assign and_tmp_40 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2])
      & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_297_nl);
  assign mux_299_nl = MUX_s_1_2_2(nor_1213_cse, and_2743_cse, MAC_LOOP_mux_11_tmp[3]);
  assign and_tmp_41 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2])
      & (MAC_LOOP_mux_11_tmp[4]) & (mux_299_nl);
  assign nor_1159_cse = ~((MAC_LOOP_mux_11_tmp[4:3]!=2'b00));
  assign and_2792_cse = (MAC_LOOP_mux_11_tmp[4:3]==2'b11);
  assign mux_301_nl = MUX_s_1_2_2(nor_1159_cse, and_2792_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_42 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[5])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_301_nl);
  assign nor_1156_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[5])
      | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2795_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[5])
      & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_303_nl = MUX_s_1_2_2((nor_1156_nl), (and_2795_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_43 = (MAC_LOOP_mux_11_tmp[4:3]==2'b11) & (mux_303_nl);
  assign mux_305_nl = MUX_s_1_2_2(nor_1159_cse, and_2792_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_44 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[5])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_305_nl);
  assign nor_1149_cse = ~((MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[5]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2801_cse = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_307_nl = MUX_s_1_2_2(nor_1149_cse, and_2801_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_45 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4])
      & (mux_307_nl);
  assign nor_1146_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[4]));
  assign and_2804_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4]);
  assign mux_309_nl = MUX_s_1_2_2((nor_1146_nl), (and_2804_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_46 = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6])
      & (mux_309_nl);
  assign mux_311_nl = MUX_s_1_2_2(nor_1149_cse, and_2801_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_47 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4])
      & (mux_311_nl);
  assign mux_313_nl = MUX_s_1_2_2(nor_1159_cse, and_2792_cse, MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_48 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[5])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_313_nl);
  assign mux_315_nl = MUX_s_1_2_2(nor_1213_cse, and_2743_cse, MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_49 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[4]) & (mux_315_nl);
  assign nor_1132_cse = ~((MAC_LOOP_mux_11_tmp[4:2]!=3'b000));
  assign and_2816_cse = (MAC_LOOP_mux_11_tmp[4:2]==3'b111);
  assign mux_317_nl = MUX_s_1_2_2(nor_1132_cse, and_2816_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_50 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6])
      & (mux_317_nl);
  assign nor_1128_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[5]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2819_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_319_nl = MUX_s_1_2_2((nor_1128_nl), (and_2819_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_51 = (MAC_LOOP_mux_11_tmp[4:2]==3'b111) & (mux_319_nl);
  assign mux_321_nl = MUX_s_1_2_2(nor_1132_cse, and_2816_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_52 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6])
      & (mux_321_nl);
  assign mux_323_nl = MUX_s_1_2_2(nor_1213_cse, and_2743_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_53 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[4]) & (mux_323_nl);
  assign nor_1117_nl = ~((MAC_LOOP_mux_11_tmp[4:1]!=4'b0000));
  assign and_2828_nl = (MAC_LOOP_mux_11_tmp[4:1]==4'b1111);
  assign mux_325_nl = MUX_s_1_2_2((nor_1117_nl), (and_2828_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_54 = (MAC_LOOP_mux_11_tmp[6:5]==2'b11) & (mux_325_nl);
  assign mux_327_nl = MUX_s_1_2_2(nor_1213_cse, and_2743_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_55 = (MAC_LOOP_mux_11_tmp[4:1]==4'b1111) & (mux_327_nl);
  assign mux_329_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[6])), (MAC_LOOP_mux_11_tmp[6]),
      MAC_LOOP_mux_11_tmp[5]);
  assign and_tmp_56 = (MAC_LOOP_mux_11_tmp[4:0]==5'b11111) & (mux_329_nl);
  assign mux_331_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[5])), (MAC_LOOP_mux_11_tmp[5]),
      MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_57 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_331_nl);
  assign nor_1105_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[3])
      | (MAC_LOOP_mux_11_tmp[4]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2840_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_333_nl = MUX_s_1_2_2((nor_1105_nl), (and_2840_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_58 = (MAC_LOOP_mux_11_tmp[5]) & (mux_333_nl);
  assign mux_335_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[5])), (MAC_LOOP_mux_11_tmp[5]),
      MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_59 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_335_nl);
  assign nor_1098_cse = ~((MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[4])
      | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2846_cse = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_337_nl = MUX_s_1_2_2(nor_1098_cse, and_2846_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_60 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[5]) & (mux_337_nl);
  assign nor_1093_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[5]));
  assign and_2849_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[5]);
  assign mux_339_nl = MUX_s_1_2_2((nor_1093_nl), (and_2849_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_61 = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_339_nl);
  assign mux_341_nl = MUX_s_1_2_2(nor_1098_cse, and_2846_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_62 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[5]) & (mux_341_nl);
  assign mux_343_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[5])), (MAC_LOOP_mux_11_tmp[5]),
      MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_63 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_343_nl);
  assign nor_1082_cse = ~((MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[4]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2858_cse = (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_345_nl = MUX_s_1_2_2(nor_1082_cse, and_2858_cse, MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_64 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[5])
      & (mux_345_nl);
  assign nor_1077_cse = ~((MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[5]));
  assign and_2861_cse = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[5]);
  assign mux_347_nl = MUX_s_1_2_2(nor_1077_cse, and_2861_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_65 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_347_nl);
  assign nor_1073_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[4])
      | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2864_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_349_nl = MUX_s_1_2_2((nor_1073_nl), (and_2864_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_66 = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[5]) & (mux_349_nl);
  assign mux_351_nl = MUX_s_1_2_2(nor_1077_cse, and_2861_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_67 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_351_nl);
  assign mux_353_nl = MUX_s_1_2_2(nor_1082_cse, and_2858_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_68 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[5])
      & (mux_353_nl);
  assign nor_1062_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[5]));
  assign and_2873_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[5]);
  assign mux_355_nl = MUX_s_1_2_2((nor_1062_nl), (and_2873_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_69 = (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6])
      & (mux_355_nl);
  assign mux_357_nl = MUX_s_1_2_2(nor_1082_cse, and_2858_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_70 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[5])
      & (mux_357_nl);
  assign mux_359_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[5])), (MAC_LOOP_mux_11_tmp[5]),
      MAC_LOOP_mux_11_tmp[3]);
  assign and_tmp_71 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2])
      & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_359_nl);
  assign nor_1052_cse = ~((MAC_LOOP_mux_11_tmp[4]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2882_cse = (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_361_nl = MUX_s_1_2_2(nor_1052_cse, and_2882_cse, MAC_LOOP_mux_11_tmp[3]);
  assign and_tmp_72 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2])
      & (MAC_LOOP_mux_11_tmp[5]) & (mux_361_nl);
  assign nor_1048_cse = ~((MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[5]));
  assign and_2885_cse = (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5]);
  assign mux_363_nl = MUX_s_1_2_2(nor_1048_cse, and_2885_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_73 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_363_nl);
  assign nor_1044_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[4])
      | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2888_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_365_nl = MUX_s_1_2_2((nor_1044_nl), (and_2888_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_74 = (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5]) & (mux_365_nl);
  assign mux_367_nl = MUX_s_1_2_2(nor_1048_cse, and_2885_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_75 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_367_nl);
  assign nor_1037_cse = ~((MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[4]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2894_cse = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_369_nl = MUX_s_1_2_2(nor_1037_cse, and_2894_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_76 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5])
      & (mux_369_nl);
  assign nor_1033_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[5]));
  assign and_2897_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5]);
  assign mux_371_nl = MUX_s_1_2_2((nor_1033_nl), (and_2897_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_77 = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6])
      & (mux_371_nl);
  assign mux_373_nl = MUX_s_1_2_2(nor_1037_cse, and_2894_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_78 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5])
      & (mux_373_nl);
  assign mux_375_nl = MUX_s_1_2_2(nor_1048_cse, and_2885_cse, MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_79 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_375_nl);
  assign mux_377_nl = MUX_s_1_2_2(nor_1052_cse, and_2882_cse, MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_80 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[5]) & (mux_377_nl);
  assign nor_1017_cse = ~((MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[5]));
  assign and_2909_cse = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5]);
  assign mux_379_nl = MUX_s_1_2_2(nor_1017_cse, and_2909_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_81 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6])
      & (mux_379_nl);
  assign nor_1012_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[4]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2912_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_381_nl = MUX_s_1_2_2((nor_1012_nl), (and_2912_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_82 = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5])
      & (mux_381_nl);
  assign mux_383_nl = MUX_s_1_2_2(nor_1017_cse, and_2909_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_83 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6])
      & (mux_383_nl);
  assign mux_385_nl = MUX_s_1_2_2(nor_1052_cse, and_2882_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_84 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[5]) & (mux_385_nl);
  assign nor_1000_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[3])
      | (MAC_LOOP_mux_11_tmp[5]));
  assign and_2921_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[5]);
  assign mux_387_nl = MUX_s_1_2_2((nor_1000_nl), (and_2921_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_85 = (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_387_nl);
  assign mux_389_nl = MUX_s_1_2_2(nor_1052_cse, and_2882_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_86 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[5]) & (mux_389_nl);
  assign mux_391_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[5])), (MAC_LOOP_mux_11_tmp[5]),
      MAC_LOOP_mux_11_tmp[4]);
  assign and_tmp_87 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2])
      & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_391_nl);
  assign mux_393_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[6])), (MAC_LOOP_mux_11_tmp[6]),
      MAC_LOOP_mux_11_tmp[4]);
  assign and_tmp_88 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2])
      & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5]) & (mux_393_nl);
  assign nor_986_cse = ~((MAC_LOOP_mux_11_tmp[5:4]!=2'b00));
  assign and_2933_cse = (MAC_LOOP_mux_11_tmp[5:4]==2'b11);
  assign mux_395_nl = MUX_s_1_2_2(nor_986_cse, and_2933_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_89 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_395_nl);
  assign nor_982_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[3])
      | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2936_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_397_nl = MUX_s_1_2_2((nor_982_nl), (and_2936_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_90 = (MAC_LOOP_mux_11_tmp[5:4]==2'b11) & (mux_397_nl);
  assign mux_399_nl = MUX_s_1_2_2(nor_986_cse, and_2933_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_91 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_399_nl);
  assign nor_975_cse = ~((MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2942_cse = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_401_nl = MUX_s_1_2_2(nor_975_cse, and_2942_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_92 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5])
      & (mux_401_nl);
  assign nor_971_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[4]) | (MAC_LOOP_mux_11_tmp[5]));
  assign and_2945_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5]);
  assign mux_403_nl = MUX_s_1_2_2((nor_971_nl), (and_2945_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_93 = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[6])
      & (mux_403_nl);
  assign mux_405_nl = MUX_s_1_2_2(nor_975_cse, and_2942_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_94 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5])
      & (mux_405_nl);
  assign mux_407_nl = MUX_s_1_2_2(nor_986_cse, and_2933_cse, MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_95 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_407_nl);
  assign nor_960_cse = ~((MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2954_cse = (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_409_nl = MUX_s_1_2_2(nor_960_cse, and_2954_cse, MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_96 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[5]) & (mux_409_nl);
  assign nor_956_cse = ~((MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[4]) | (MAC_LOOP_mux_11_tmp[5]));
  assign and_2957_cse = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5]);
  assign mux_411_nl = MUX_s_1_2_2(nor_956_cse, and_2957_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_97 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[6])
      & (mux_411_nl);
  assign nor_952_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2960_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_413_nl = MUX_s_1_2_2((nor_952_nl), (and_2960_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_98 = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5])
      & (mux_413_nl);
  assign mux_415_nl = MUX_s_1_2_2(nor_956_cse, and_2957_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_99 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[6])
      & (mux_415_nl);
  assign mux_417_nl = MUX_s_1_2_2(nor_960_cse, and_2954_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_100 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[5]) & (mux_417_nl);
  assign nor_943_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[4])
      | (MAC_LOOP_mux_11_tmp[5]));
  assign and_2969_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[5]);
  assign mux_419_nl = MUX_s_1_2_2((nor_943_nl), (and_2969_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_101 = (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_419_nl);
  assign mux_421_nl = MUX_s_1_2_2(nor_960_cse, and_2954_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_102 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[5]) & (mux_421_nl);
  assign mux_423_nl = MUX_s_1_2_2(nor_986_cse, and_2933_cse, MAC_LOOP_mux_11_tmp[3]);
  assign and_tmp_103 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2])
      & (MAC_LOOP_mux_11_tmp[6]) & (mux_423_nl);
  assign mux_425_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[6])), (MAC_LOOP_mux_11_tmp[6]),
      MAC_LOOP_mux_11_tmp[3]);
  assign and_tmp_104 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2])
      & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5]) & (mux_425_nl);
  assign nor_931_cse = ~((MAC_LOOP_mux_11_tmp[5:3]!=3'b000));
  assign and_2981_cse = (MAC_LOOP_mux_11_tmp[5:3]==3'b111);
  assign mux_427_nl = MUX_s_1_2_2(nor_931_cse, and_2981_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_105 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[6])
      & (mux_427_nl);
  assign nor_927_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2984_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_429_nl = MUX_s_1_2_2((nor_927_nl), (and_2984_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_106 = (MAC_LOOP_mux_11_tmp[5:3]==3'b111) & (mux_429_nl);
  assign mux_431_nl = MUX_s_1_2_2(nor_931_cse, and_2981_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_107 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[6])
      & (mux_431_nl);
  assign nor_921_cse = ~((MAC_LOOP_mux_11_tmp[2]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_2990_cse = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_433_nl = MUX_s_1_2_2(nor_921_cse, and_2990_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_108 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[5]) & (mux_433_nl);
  assign nor_918_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[3]) | (MAC_LOOP_mux_11_tmp[4])
      | (MAC_LOOP_mux_11_tmp[5]));
  assign and_2993_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[5]);
  assign mux_435_nl = MUX_s_1_2_2((nor_918_nl), (and_2993_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_109 = (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_435_nl);
  assign mux_437_nl = MUX_s_1_2_2(nor_921_cse, and_2990_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_110 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4])
      & (MAC_LOOP_mux_11_tmp[5]) & (mux_437_nl);
  assign mux_439_nl = MUX_s_1_2_2(nor_931_cse, and_2981_cse, MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_111 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[6])
      & (mux_439_nl);
  assign mux_441_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[6])), (MAC_LOOP_mux_11_tmp[6]),
      MAC_LOOP_mux_11_tmp[2]);
  assign and_tmp_112 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5]) & (mux_441_nl);
  assign nor_905_cse = ~((MAC_LOOP_mux_11_tmp[5:2]!=4'b0000));
  assign and_3005_cse = (MAC_LOOP_mux_11_tmp[5:2]==4'b1111);
  assign mux_443_nl = MUX_s_1_2_2(nor_905_cse, and_3005_cse, MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_113 = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_443_nl);
  assign nor_900_nl = ~((MAC_LOOP_mux_11_tmp[1]) | (MAC_LOOP_mux_11_tmp[6]));
  assign and_3008_nl = (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[6]);
  assign mux_445_nl = MUX_s_1_2_2((nor_900_nl), (and_3008_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_114 = (MAC_LOOP_mux_11_tmp[5:2]==4'b1111) & (mux_445_nl);
  assign mux_447_nl = MUX_s_1_2_2(nor_905_cse, and_3005_cse, MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_115 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_447_nl);
  assign mux_449_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[6])), (MAC_LOOP_mux_11_tmp[6]),
      MAC_LOOP_mux_11_tmp[1]);
  assign and_tmp_116 = (MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
      & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5]) & (mux_449_nl);
  assign nor_891_nl = ~((MAC_LOOP_mux_11_tmp[5:1]!=5'b00000));
  assign and_3016_nl = (MAC_LOOP_mux_11_tmp[5:1]==5'b11111);
  assign mux_451_nl = MUX_s_1_2_2((nor_891_nl), (and_3016_nl), MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_117 = (MAC_LOOP_mux_11_tmp[6]) & (mux_451_nl);
  assign mux_453_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[6])), (MAC_LOOP_mux_11_tmp[6]),
      MAC_LOOP_mux_11_tmp[0]);
  assign and_tmp_118 = (MAC_LOOP_mux_11_tmp[5:1]==5'b11111) & (mux_453_nl);
  always @(posedge clk) begin
    if ( rst ) begin
      y_rsci_idat_0 <= 1'b0;
    end
    else if ( fsm_output[3] ) begin
      y_rsci_idat_0 <= (z_out_2[0]) | nor_ovfl_sva_1 | and_unfl_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      y_rsci_idat_7_1 <= 7'b0000000;
    end
    else if ( fsm_output[3] ) begin
      y_rsci_idat_7_1 <= ~(MUX_v_7_2_2((nor_5_nl), 7'b1111111, and_unfl_sva_1));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      y_rsci_idat_8 <= 1'b0;
    end
    else if ( fsm_output[3] ) begin
      y_rsci_idat_8 <= z_out_2[14];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_sample_sva <= 3'b000;
    end
    else if ( ~((fsm_output[2:1]!=2'b00)) ) begin
      i_sample_sva <= i_sample_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_126_lpi_2 <= 3'b000;
    end
    else if ( (~(((MAC_LOOP_mux_11_tmp[6:1]==6'b111111)) | ((acc_2_tmp_7_1[6:1]==6'b111111))))
        & (~ (fsm_output[2])) & (MAC_LOOP_n_6_0_sva==7'b1111110) ) begin
      x_126_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_125_lpi_2 <= 3'b000;
    end
    else if ( (~(((MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[3])
        & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]))
        | (((acc_2_tmp_7_1[1:0]!=2'b00)) & (acc_2_tmp_7_1[6:2]==5'b11111)))) & (fsm_output[1])
        & (MAC_LOOP_n_6_0_sva==7'b1111101) ) begin
      x_125_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_1_lpi_2 <= 3'b000;
    end
    else if ( (mux_221_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & nor_1309_cse & (~ (MAC_LOOP_n_6_0_sva[5])) & (MAC_LOOP_n_6_0_sva[0]) )
        begin
      x_1_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_124_lpi_2 <= 3'b000;
    end
    else if ( (~((((acc_2_tmp_7_1[1:0]!=2'b01)) & (acc_2_tmp_7_1[6:2]==5'b11111))
        | ((MAC_LOOP_mux_11_tmp[6:2]==5'b11111) & (mux_222_nl)))) & (fsm_output[1])
        & (MAC_LOOP_n_6_0_sva==7'b1111100) ) begin
      x_124_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_2_lpi_2 <= 3'b000;
    end
    else if ( (mux_224_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & nor_1309_cse & nor_1303_cse ) begin
      x_2_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_123_lpi_2 <= 3'b000;
    end
    else if ( (~(((MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3])
        & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]))
        | (((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[0])) & (acc_2_tmp_7_1[5]) & (acc_2_tmp_7_1[6])
        & (acc_2_tmp_7_1[3]) & (acc_2_tmp_7_1[4]) & (acc_2_tmp_7_1[1])))) & (fsm_output[1])
        & (MAC_LOOP_n_6_0_sva==7'b1111011) ) begin
      x_123_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_3_lpi_2 <= 3'b000;
    end
    else if ( (mux_226_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & nor_1309_cse & (~ (MAC_LOOP_n_6_0_sva[5])) & (MAC_LOOP_n_6_0_sva[0]) )
        begin
      x_3_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_122_lpi_2 <= 3'b000;
    end
    else if ( (~((((acc_2_tmp_7_1[2]) | (~ (acc_2_tmp_7_1[0]))) & (acc_2_tmp_7_1[5])
        & (acc_2_tmp_7_1[6]) & (acc_2_tmp_7_1[3]) & (acc_2_tmp_7_1[4]) & (acc_2_tmp_7_1[1]))
        | ((MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4])
        & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_227_nl)))) &
        (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1111010) ) begin
      x_122_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_4_lpi_2 <= 3'b000;
    end
    else if ( (mux_229_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b010)
        & nor_1309_cse & nor_1303_cse ) begin
      x_4_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_121_lpi_2 <= 3'b000;
    end
    else if ( (mux_231_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1111001) )
        begin
      x_121_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_5_lpi_2 <= 3'b000;
    end
    else if ( (mux_233_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b010)
        & nor_1309_cse & (~ (MAC_LOOP_n_6_0_sva[5])) & (MAC_LOOP_n_6_0_sva[0]) )
        begin
      x_5_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_120_lpi_2 <= 3'b000;
    end
    else if ( (mux_235_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1111000) )
        begin
      x_120_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_6_lpi_2 <= 3'b000;
    end
    else if ( (mux_237_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b011)
        & nor_1309_cse & nor_1303_cse ) begin
      x_6_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_119_lpi_2 <= 3'b000;
    end
    else if ( (~(((MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2])
        & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]))
        | (((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[0])) & (acc_2_tmp_7_1[5]) & (acc_2_tmp_7_1[6])
        & (acc_2_tmp_7_1[4]) & (acc_2_tmp_7_1[2]) & (acc_2_tmp_7_1[1])))) & (fsm_output[1])
        & (MAC_LOOP_n_6_0_sva==7'b1110111) ) begin
      x_119_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_7_lpi_2 <= 3'b000;
    end
    else if ( (mux_239_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b011)
        & nor_1309_cse & (~ (MAC_LOOP_n_6_0_sva[5])) & (MAC_LOOP_n_6_0_sva[0]) )
        begin
      x_7_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_118_lpi_2 <= 3'b000;
    end
    else if ( (~((((acc_2_tmp_7_1[3]) | (~ (acc_2_tmp_7_1[0]))) & (acc_2_tmp_7_1[5])
        & (acc_2_tmp_7_1[6]) & (acc_2_tmp_7_1[4]) & (acc_2_tmp_7_1[2]) & (acc_2_tmp_7_1[1]))
        | ((MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2]) & (MAC_LOOP_mux_11_tmp[4])
        & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]) & (mux_240_nl)))) &
        (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1110110) ) begin
      x_118_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_8_lpi_2 <= 3'b000;
    end
    else if ( (mux_242_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b100)
        & nor_1309_cse & nor_1303_cse ) begin
      x_8_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_117_lpi_2 <= 3'b000;
    end
    else if ( (mux_244_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1110101) )
        begin
      x_117_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_9_lpi_2 <= 3'b000;
    end
    else if ( (mux_246_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b100)
        & nor_1309_cse & (~ (MAC_LOOP_n_6_0_sva[5])) & (MAC_LOOP_n_6_0_sva[0]) )
        begin
      x_9_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_116_lpi_2 <= 3'b000;
    end
    else if ( (mux_248_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1110100) )
        begin
      x_116_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_10_lpi_2 <= 3'b000;
    end
    else if ( (mux_250_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b101)
        & nor_1309_cse & nor_1303_cse ) begin
      x_10_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_115_lpi_2 <= 3'b000;
    end
    else if ( (mux_252_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (MAC_LOOP_n_6_0_sva[6]) & (MAC_LOOP_n_6_0_sva[5])
        & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_115_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_11_lpi_2 <= 3'b000;
    end
    else if ( (mux_254_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b101)
        & nor_1309_cse & (~ (MAC_LOOP_n_6_0_sva[5])) & (MAC_LOOP_n_6_0_sva[0]) )
        begin
      x_11_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_114_lpi_2 <= 3'b000;
    end
    else if ( (mux_256_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (MAC_LOOP_n_6_0_sva[6]) & (MAC_LOOP_n_6_0_sva[5])
        & (~ (MAC_LOOP_n_6_0_sva[0])) ) begin
      x_114_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_12_lpi_2 <= 3'b000;
    end
    else if ( (mux_258_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b110)
        & nor_1309_cse & nor_1303_cse ) begin
      x_12_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_113_lpi_2 <= 3'b000;
    end
    else if ( (mux_260_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (MAC_LOOP_n_6_0_sva[6]) & (MAC_LOOP_n_6_0_sva[5])
        & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_113_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_13_lpi_2 <= 3'b000;
    end
    else if ( (mux_262_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b110)
        & nor_1309_cse & (~ (MAC_LOOP_n_6_0_sva[5])) & (MAC_LOOP_n_6_0_sva[0]) )
        begin
      x_13_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_112_lpi_2 <= 3'b000;
    end
    else if ( (mux_264_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (MAC_LOOP_n_6_0_sva[6]) & (MAC_LOOP_n_6_0_sva[5])
        & (~ (MAC_LOOP_n_6_0_sva[0])) ) begin
      x_112_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_14_lpi_2 <= 3'b000;
    end
    else if ( (mux_266_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b111)
        & nor_1309_cse & nor_1303_cse ) begin
      x_14_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_111_lpi_2 <= 3'b000;
    end
    else if ( (~(((MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2])
        & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[5]) & (MAC_LOOP_mux_11_tmp[6]))
        | (((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[0])) & (acc_2_tmp_7_1[5]) & (acc_2_tmp_7_1[6])
        & (acc_2_tmp_7_1[2]) & (acc_2_tmp_7_1[3]) & (acc_2_tmp_7_1[1])))) & (fsm_output[1])
        & (MAC_LOOP_n_6_0_sva==7'b1101111) ) begin
      x_111_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_15_lpi_2 <= 3'b000;
    end
    else if ( (mux_268_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b111)
        & nor_1309_cse & (~ (MAC_LOOP_n_6_0_sva[5])) & (MAC_LOOP_n_6_0_sva[0]) )
        begin
      x_15_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_110_lpi_2 <= 3'b000;
    end
    else if ( (~ (mux_270_nl)) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1101110)
        ) begin
      x_110_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_16_lpi_2 <= 3'b000;
    end
    else if ( (mux_272_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (~ (MAC_LOOP_n_6_0_sva[6])) & nor_1303_cse )
        begin
      x_16_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_109_lpi_2 <= 3'b000;
    end
    else if ( (mux_274_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1101101) )
        begin
      x_109_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_17_lpi_2 <= 3'b000;
    end
    else if ( (mux_276_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (~ (MAC_LOOP_n_6_0_sva[6])) & (~ (MAC_LOOP_n_6_0_sva[5]))
        & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_17_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_108_lpi_2 <= 3'b000;
    end
    else if ( (mux_278_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1101100) )
        begin
      x_108_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_18_lpi_2 <= 3'b000;
    end
    else if ( (mux_280_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (~ (MAC_LOOP_n_6_0_sva[6])) & nor_1303_cse )
        begin
      x_18_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_107_lpi_2 <= 3'b000;
    end
    else if ( (mux_282_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1101011) )
        begin
      x_107_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_19_lpi_2 <= 3'b000;
    end
    else if ( (mux_284_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (~ (MAC_LOOP_n_6_0_sva[6])) & (~ (MAC_LOOP_n_6_0_sva[5]))
        & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_19_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_106_lpi_2 <= 3'b000;
    end
    else if ( (mux_286_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1101010) )
        begin
      x_106_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_20_lpi_2 <= 3'b000;
    end
    else if ( (mux_288_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & (MAC_LOOP_n_6_0_sva[2])
        & (~ (MAC_LOOP_n_6_0_sva[3])) & (MAC_LOOP_n_6_0_sva[4]) & (~ (MAC_LOOP_n_6_0_sva[6]))
        & nor_1303_cse ) begin
      x_20_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_105_lpi_2 <= 3'b000;
    end
    else if ( (mux_290_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1101001) )
        begin
      x_105_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_21_lpi_2 <= 3'b000;
    end
    else if ( (mux_292_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0010101) )
        begin
      x_21_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_104_lpi_2 <= 3'b000;
    end
    else if ( (mux_294_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1101000) )
        begin
      x_104_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_22_lpi_2 <= 3'b000;
    end
    else if ( (mux_296_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & (MAC_LOOP_n_6_0_sva[2])
        & (~ (MAC_LOOP_n_6_0_sva[3])) & (MAC_LOOP_n_6_0_sva[4]) & (~ (MAC_LOOP_n_6_0_sva[6]))
        & nor_1303_cse ) begin
      x_22_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_103_lpi_2 <= 3'b000;
    end
    else if ( (mux_298_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1100111) )
        begin
      x_103_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_23_lpi_2 <= 3'b000;
    end
    else if ( (mux_300_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0010111) )
        begin
      x_23_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_102_lpi_2 <= 3'b000;
    end
    else if ( (mux_302_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1100110) )
        begin
      x_102_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_24_lpi_2 <= 3'b000;
    end
    else if ( (mux_304_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & (~ (MAC_LOOP_n_6_0_sva[2]))
        & (MAC_LOOP_n_6_0_sva[3]) & (MAC_LOOP_n_6_0_sva[4]) & (~ (MAC_LOOP_n_6_0_sva[6]))
        & nor_1303_cse ) begin
      x_24_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_101_lpi_2 <= 3'b000;
    end
    else if ( (mux_306_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1100101) )
        begin
      x_101_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_25_lpi_2 <= 3'b000;
    end
    else if ( (mux_308_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0011001) )
        begin
      x_25_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_100_lpi_2 <= 3'b000;
    end
    else if ( (mux_310_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1100100) )
        begin
      x_100_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_26_lpi_2 <= 3'b000;
    end
    else if ( (mux_312_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & (~ (MAC_LOOP_n_6_0_sva[2]))
        & (MAC_LOOP_n_6_0_sva[3]) & (MAC_LOOP_n_6_0_sva[4]) & (~ (MAC_LOOP_n_6_0_sva[6]))
        & nor_1303_cse ) begin
      x_26_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_99_lpi_2 <= 3'b000;
    end
    else if ( (mux_314_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & (~ (MAC_LOOP_n_6_0_sva[4])) & (MAC_LOOP_n_6_0_sva[6]) & (MAC_LOOP_n_6_0_sva[5])
        & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_99_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_27_lpi_2 <= 3'b000;
    end
    else if ( (mux_316_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0011011) )
        begin
      x_27_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_98_lpi_2 <= 3'b000;
    end
    else if ( (mux_318_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & (~ (MAC_LOOP_n_6_0_sva[4])) & (MAC_LOOP_n_6_0_sva[6]) & (MAC_LOOP_n_6_0_sva[5])
        & (~ (MAC_LOOP_n_6_0_sva[0])) ) begin
      x_98_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_28_lpi_2 <= 3'b000;
    end
    else if ( (mux_320_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & (MAC_LOOP_n_6_0_sva[2])
        & (MAC_LOOP_n_6_0_sva[3]) & (MAC_LOOP_n_6_0_sva[4]) & (~ (MAC_LOOP_n_6_0_sva[6]))
        & nor_1303_cse ) begin
      x_28_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_97_lpi_2 <= 3'b000;
    end
    else if ( (mux_322_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & (~ (MAC_LOOP_n_6_0_sva[4])) & (MAC_LOOP_n_6_0_sva[6]) & (MAC_LOOP_n_6_0_sva[5])
        & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_97_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_29_lpi_2 <= 3'b000;
    end
    else if ( (mux_324_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0011101) )
        begin
      x_29_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_96_lpi_2 <= 3'b000;
    end
    else if ( (mux_326_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & (~ (MAC_LOOP_n_6_0_sva[4])) & (MAC_LOOP_n_6_0_sva[6]) & (MAC_LOOP_n_6_0_sva[5])
        & (~ (MAC_LOOP_n_6_0_sva[0])) ) begin
      x_96_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_30_lpi_2 <= 3'b000;
    end
    else if ( (mux_328_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & (MAC_LOOP_n_6_0_sva[2])
        & (MAC_LOOP_n_6_0_sva[3]) & (MAC_LOOP_n_6_0_sva[4]) & (~ (MAC_LOOP_n_6_0_sva[6]))
        & nor_1303_cse ) begin
      x_30_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_95_lpi_2 <= 3'b000;
    end
    else if ( (~(((MAC_LOOP_mux_11_tmp[0]) & (MAC_LOOP_mux_11_tmp[1]) & (MAC_LOOP_mux_11_tmp[2])
        & (MAC_LOOP_mux_11_tmp[3]) & (MAC_LOOP_mux_11_tmp[4]) & (MAC_LOOP_mux_11_tmp[6]))
        | (((acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[0])) & (acc_2_tmp_7_1[6]) & (acc_2_tmp_7_1[4])
        & (acc_2_tmp_7_1[2]) & (acc_2_tmp_7_1[3]) & (acc_2_tmp_7_1[1])))) & (fsm_output[1])
        & (MAC_LOOP_n_6_0_sva==7'b1011111) ) begin
      x_95_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_31_lpi_2 <= 3'b000;
    end
    else if ( (mux_330_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0011111) )
        begin
      x_31_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_94_lpi_2 <= 3'b000;
    end
    else if ( (~ (mux_332_nl)) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & (MAC_LOOP_n_6_0_sva[2])
        & (MAC_LOOP_n_6_0_sva[3]) & (MAC_LOOP_n_6_0_sva[4]) & (MAC_LOOP_n_6_0_sva[6])
        & nor_1303_cse ) begin
      x_94_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_32_lpi_2 <= 3'b000;
    end
    else if ( (mux_334_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (~ (MAC_LOOP_n_6_0_sva[0])) )
        begin
      x_32_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_93_lpi_2 <= 3'b000;
    end
    else if ( (mux_336_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1011101) )
        begin
      x_93_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_33_lpi_2 <= 3'b000;
    end
    else if ( (mux_338_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_33_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_92_lpi_2 <= 3'b000;
    end
    else if ( (mux_340_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & (MAC_LOOP_n_6_0_sva[2])
        & (MAC_LOOP_n_6_0_sva[3]) & (MAC_LOOP_n_6_0_sva[4]) & (MAC_LOOP_n_6_0_sva[6])
        & nor_1303_cse ) begin
      x_92_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_34_lpi_2 <= 3'b000;
    end
    else if ( (mux_342_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (~ (MAC_LOOP_n_6_0_sva[0])) )
        begin
      x_34_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_91_lpi_2 <= 3'b000;
    end
    else if ( (mux_344_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1011011) )
        begin
      x_91_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_35_lpi_2 <= 3'b000;
    end
    else if ( (mux_346_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_35_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_90_lpi_2 <= 3'b000;
    end
    else if ( (mux_348_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & (~ (MAC_LOOP_n_6_0_sva[2]))
        & (MAC_LOOP_n_6_0_sva[3]) & (MAC_LOOP_n_6_0_sva[4]) & (MAC_LOOP_n_6_0_sva[6])
        & nor_1303_cse ) begin
      x_90_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_36_lpi_2 <= 3'b000;
    end
    else if ( (mux_350_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b010)
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (~ (MAC_LOOP_n_6_0_sva[0])) )
        begin
      x_36_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_89_lpi_2 <= 3'b000;
    end
    else if ( (mux_352_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1011001) )
        begin
      x_89_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_37_lpi_2 <= 3'b000;
    end
    else if ( (mux_354_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b010)
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_37_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_88_lpi_2 <= 3'b000;
    end
    else if ( (mux_356_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & (~ (MAC_LOOP_n_6_0_sva[2]))
        & (MAC_LOOP_n_6_0_sva[3]) & (MAC_LOOP_n_6_0_sva[4]) & (MAC_LOOP_n_6_0_sva[6])
        & nor_1303_cse ) begin
      x_88_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_38_lpi_2 <= 3'b000;
    end
    else if ( (mux_358_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b011)
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (~ (MAC_LOOP_n_6_0_sva[0])) )
        begin
      x_38_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_87_lpi_2 <= 3'b000;
    end
    else if ( (mux_360_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1010111) )
        begin
      x_87_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_39_lpi_2 <= 3'b000;
    end
    else if ( (mux_362_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b011)
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_39_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_86_lpi_2 <= 3'b000;
    end
    else if ( (mux_364_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & (MAC_LOOP_n_6_0_sva[2])
        & (~ (MAC_LOOP_n_6_0_sva[3])) & (MAC_LOOP_n_6_0_sva[4]) & (MAC_LOOP_n_6_0_sva[6])
        & nor_1303_cse ) begin
      x_86_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_40_lpi_2 <= 3'b000;
    end
    else if ( (mux_366_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b100)
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (~ (MAC_LOOP_n_6_0_sva[0])) )
        begin
      x_40_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_85_lpi_2 <= 3'b000;
    end
    else if ( (mux_368_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1010101) )
        begin
      x_85_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_41_lpi_2 <= 3'b000;
    end
    else if ( (mux_370_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b100)
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_41_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_84_lpi_2 <= 3'b000;
    end
    else if ( (mux_372_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & (MAC_LOOP_n_6_0_sva[2])
        & (~ (MAC_LOOP_n_6_0_sva[3])) & (MAC_LOOP_n_6_0_sva[4]) & (MAC_LOOP_n_6_0_sva[6])
        & nor_1303_cse ) begin
      x_84_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_42_lpi_2 <= 3'b000;
    end
    else if ( (mux_374_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b101)
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (~ (MAC_LOOP_n_6_0_sva[0])) )
        begin
      x_42_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_83_lpi_2 <= 3'b000;
    end
    else if ( (mux_376_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (MAC_LOOP_n_6_0_sva[6]) & (~ (MAC_LOOP_n_6_0_sva[5]))
        & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_83_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_43_lpi_2 <= 3'b000;
    end
    else if ( (mux_378_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b101)
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_43_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_82_lpi_2 <= 3'b000;
    end
    else if ( (mux_380_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (MAC_LOOP_n_6_0_sva[6]) & nor_1303_cse ) begin
      x_82_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_44_lpi_2 <= 3'b000;
    end
    else if ( (mux_382_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b110)
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (~ (MAC_LOOP_n_6_0_sva[0])) )
        begin
      x_44_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_81_lpi_2 <= 3'b000;
    end
    else if ( (mux_384_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (MAC_LOOP_n_6_0_sva[6]) & (~ (MAC_LOOP_n_6_0_sva[5]))
        & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_81_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_45_lpi_2 <= 3'b000;
    end
    else if ( (mux_386_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b110)
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_45_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_80_lpi_2 <= 3'b000;
    end
    else if ( (mux_388_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (MAC_LOOP_n_6_0_sva[6]) & nor_1303_cse ) begin
      x_80_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_46_lpi_2 <= 3'b000;
    end
    else if ( (mux_390_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b111)
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (~ (MAC_LOOP_n_6_0_sva[0])) )
        begin
      x_46_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_79_lpi_2 <= 3'b000;
    end
    else if ( (mux_392_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1001111) )
        begin
      x_79_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_47_lpi_2 <= 3'b000;
    end
    else if ( (mux_394_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[3:1]==3'b111)
        & nor_1309_cse & (MAC_LOOP_n_6_0_sva[5]) & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_47_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_78_lpi_2 <= 3'b000;
    end
    else if ( (mux_396_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & (MAC_LOOP_n_6_0_sva[2])
        & (MAC_LOOP_n_6_0_sva[3]) & (~ (MAC_LOOP_n_6_0_sva[4])) & (MAC_LOOP_n_6_0_sva[6])
        & nor_1303_cse ) begin
      x_78_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_48_lpi_2 <= 3'b000;
    end
    else if ( (mux_398_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (~ (MAC_LOOP_n_6_0_sva[6])) & (MAC_LOOP_n_6_0_sva[5])
        & (~ (MAC_LOOP_n_6_0_sva[0])) ) begin
      x_48_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_77_lpi_2 <= 3'b000;
    end
    else if ( (mux_400_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1001101) )
        begin
      x_77_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_49_lpi_2 <= 3'b000;
    end
    else if ( (mux_402_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (~ (MAC_LOOP_n_6_0_sva[6])) & (MAC_LOOP_n_6_0_sva[5])
        & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_49_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_76_lpi_2 <= 3'b000;
    end
    else if ( (mux_404_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & (MAC_LOOP_n_6_0_sva[2])
        & (MAC_LOOP_n_6_0_sva[3]) & (~ (MAC_LOOP_n_6_0_sva[4])) & (MAC_LOOP_n_6_0_sva[6])
        & nor_1303_cse ) begin
      x_76_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_50_lpi_2 <= 3'b000;
    end
    else if ( (mux_406_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (~ (MAC_LOOP_n_6_0_sva[6])) & (MAC_LOOP_n_6_0_sva[5])
        & (~ (MAC_LOOP_n_6_0_sva[0])) ) begin
      x_50_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_75_lpi_2 <= 3'b000;
    end
    else if ( (mux_408_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1001011) )
        begin
      x_75_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_51_lpi_2 <= 3'b000;
    end
    else if ( (mux_410_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & (MAC_LOOP_n_6_0_sva[4]) & (~ (MAC_LOOP_n_6_0_sva[6])) & (MAC_LOOP_n_6_0_sva[5])
        & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_51_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_74_lpi_2 <= 3'b000;
    end
    else if ( (mux_412_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & (~ (MAC_LOOP_n_6_0_sva[2]))
        & (MAC_LOOP_n_6_0_sva[3]) & (~ (MAC_LOOP_n_6_0_sva[4])) & (MAC_LOOP_n_6_0_sva[6])
        & nor_1303_cse ) begin
      x_74_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_52_lpi_2 <= 3'b000;
    end
    else if ( (mux_414_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0110100) )
        begin
      x_52_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_73_lpi_2 <= 3'b000;
    end
    else if ( (mux_416_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1001001) )
        begin
      x_73_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_53_lpi_2 <= 3'b000;
    end
    else if ( (mux_418_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0110101) )
        begin
      x_53_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_72_lpi_2 <= 3'b000;
    end
    else if ( (mux_420_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & (~ (MAC_LOOP_n_6_0_sva[2]))
        & (MAC_LOOP_n_6_0_sva[3]) & (~ (MAC_LOOP_n_6_0_sva[4])) & (MAC_LOOP_n_6_0_sva[6])
        & nor_1303_cse ) begin
      x_72_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_54_lpi_2 <= 3'b000;
    end
    else if ( (mux_422_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0110110) )
        begin
      x_54_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_71_lpi_2 <= 3'b000;
    end
    else if ( (mux_424_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1000111) )
        begin
      x_71_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_55_lpi_2 <= 3'b000;
    end
    else if ( (mux_426_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0110111) )
        begin
      x_55_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_70_lpi_2 <= 3'b000;
    end
    else if ( (mux_428_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & (MAC_LOOP_n_6_0_sva[2])
        & (~ (MAC_LOOP_n_6_0_sva[3])) & (~ (MAC_LOOP_n_6_0_sva[4])) & (MAC_LOOP_n_6_0_sva[6])
        & nor_1303_cse ) begin
      x_70_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_56_lpi_2 <= 3'b000;
    end
    else if ( (mux_430_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0111000) )
        begin
      x_56_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_69_lpi_2 <= 3'b000;
    end
    else if ( (mux_432_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b1000101) )
        begin
      x_69_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_57_lpi_2 <= 3'b000;
    end
    else if ( (mux_434_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0111001) )
        begin
      x_57_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_68_lpi_2 <= 3'b000;
    end
    else if ( (mux_436_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & (MAC_LOOP_n_6_0_sva[2])
        & (~ (MAC_LOOP_n_6_0_sva[3])) & (~ (MAC_LOOP_n_6_0_sva[4])) & (MAC_LOOP_n_6_0_sva[6])
        & nor_1303_cse ) begin
      x_68_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_58_lpi_2 <= 3'b000;
    end
    else if ( (mux_438_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0111010) )
        begin
      x_58_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_67_lpi_2 <= 3'b000;
    end
    else if ( (mux_440_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & (~ (MAC_LOOP_n_6_0_sva[4])) & (MAC_LOOP_n_6_0_sva[6]) & (~ (MAC_LOOP_n_6_0_sva[5]))
        & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_67_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_59_lpi_2 <= 3'b000;
    end
    else if ( (mux_442_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0111011) )
        begin
      x_59_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_66_lpi_2 <= 3'b000;
    end
    else if ( (mux_444_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva[1]) & nor_1308_cse
        & (~ (MAC_LOOP_n_6_0_sva[4])) & (MAC_LOOP_n_6_0_sva[6]) & nor_1303_cse )
        begin
      x_66_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_60_lpi_2 <= 3'b000;
    end
    else if ( (mux_446_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0111100) )
        begin
      x_60_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_65_lpi_2 <= 3'b000;
    end
    else if ( (mux_448_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & (~ (MAC_LOOP_n_6_0_sva[4])) & (MAC_LOOP_n_6_0_sva[6]) & (~ (MAC_LOOP_n_6_0_sva[5]))
        & (MAC_LOOP_n_6_0_sva[0]) ) begin
      x_65_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_61_lpi_2 <= 3'b000;
    end
    else if ( (mux_450_nl) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0111101) )
        begin
      x_61_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_64_lpi_2 <= 3'b000;
    end
    else if ( (mux_452_nl) & (fsm_output[1]) & (~ (MAC_LOOP_n_6_0_sva[1])) & nor_1308_cse
        & (~ (MAC_LOOP_n_6_0_sva[4])) & (MAC_LOOP_n_6_0_sva[6]) & nor_1303_cse )
        begin
      x_64_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_62_lpi_2 <= 3'b000;
    end
    else if ( (~ (mux_454_nl)) & (fsm_output[1]) & (MAC_LOOP_n_6_0_sva==7'b0111110)
        ) begin
      x_62_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_63_lpi_2 <= 3'b000;
    end
    else if ( (~(((MAC_LOOP_mux_11_tmp[5:0]==6'b111111)) | (((acc_2_tmp_7_1[6]) |
        (acc_2_tmp_7_1[0])) & (acc_2_tmp_7_1[5:1]==5'b11111)))) & (fsm_output[1])
        & (MAC_LOOP_n_6_0_sva==7'b0111111) ) begin
      x_63_lpi_2 <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      x_0_sva <= 3'b000;
    end
    else if ( fsm_output[2] ) begin
      x_0_sva <= i_sample_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      y_rsc_triosy_obj_ld <= 1'b0;
      reg_b_rsc_triosy_obj_ld_cse <= 1'b0;
      MAC_LOOP_n_6_0_sva <= 7'b0000000;
      sum_sva <= 20'b00000000000000000000;
    end
    else begin
      y_rsc_triosy_obj_ld <= fsm_output[3];
      reg_b_rsc_triosy_obj_ld_cse <= (~ z_out_1_7) & (fsm_output[2]);
      MAC_LOOP_n_6_0_sva <= MUX_v_7_2_2(7'b0000000, (SHIFT_LOOP_n_SHIFT_LOOP_n_mux_nl),
          (MAC_LOOP_n_nor_nl));
      sum_sva <= MUX_v_20_2_2(20'b00000000000000000000, z_out_2, (fsm_output[2]));
    end
  end
  assign nor_5_nl = ~(MUX_v_7_2_2((z_out_2[7:1]), 7'b1111111, nor_ovfl_sva_1));
  assign nor_1306_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4])
      | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6]) | (~ (acc_2_tmp_7_1[0])))) | and_tmp);
  assign nor_1307_nl = ~(and_2667_cse | and_tmp);
  assign mux_221_nl = MUX_s_1_2_2((nor_1306_nl), (nor_1307_nl), acc_2_tmp_7_1[1]);
  assign mux_222_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[1])), (MAC_LOOP_mux_11_tmp[1]),
      MAC_LOOP_mux_11_tmp[0]);
  assign nor_1299_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5])
      | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[1])))) | and_tmp_2);
  assign nor_1300_nl = ~(and_2671_cse | and_tmp_2);
  assign mux_224_nl = MUX_s_1_2_2((nor_1299_nl), (nor_1300_nl), acc_2_tmp_7_1[2]);
  assign nor_1293_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5])
      | (acc_2_tmp_7_1[6]) | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[1])))) |
      and_tmp_3);
  assign nor_1294_nl = ~(and_2671_cse | and_tmp_3);
  assign mux_226_nl = MUX_s_1_2_2((nor_1293_nl), (nor_1294_nl), acc_2_tmp_7_1[2]);
  assign mux_227_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[2])), (MAC_LOOP_mux_11_tmp[2]),
      MAC_LOOP_mux_11_tmp[0]);
  assign nor_1287_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5])
      | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[2])))) | and_tmp_5);
  assign nor_1288_nl = ~(and_2667_cse | and_tmp_5);
  assign mux_229_nl = MUX_s_1_2_2((nor_1287_nl), (nor_1288_nl), acc_2_tmp_7_1[1]);
  assign nor_1285_nl = ~(((~ (acc_2_tmp_7_1[2])) & (acc_2_tmp_7_1[0]) & (acc_2_tmp_7_1[6])
      & (acc_2_tmp_7_1[5]) & (acc_2_tmp_7_1[4]) & (acc_2_tmp_7_1[3])) | and_tmp_6);
  assign nor_1286_nl = ~(and_2667_cse | and_tmp_6);
  assign mux_231_nl = MUX_s_1_2_2((nor_1285_nl), (nor_1286_nl), acc_2_tmp_7_1[1]);
  assign nor_1281_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5])
      | (acc_2_tmp_7_1[6]) | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[2])))) |
      and_tmp_7);
  assign nor_1282_nl = ~(and_2667_cse | and_tmp_7);
  assign mux_233_nl = MUX_s_1_2_2((nor_1281_nl), (nor_1282_nl), acc_2_tmp_7_1[1]);
  assign nor_1278_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[6]))
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[3]))))
      | and_tmp_8);
  assign nor_1279_nl = ~(and_2667_cse | and_tmp_8);
  assign mux_235_nl = MUX_s_1_2_2((nor_1278_nl), (nor_1279_nl), acc_2_tmp_7_1[1]);
  assign nor_1273_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[2])))) |
      and_tmp_9);
  assign nor_1274_nl = ~(and_2691_cse | and_tmp_9);
  assign mux_237_nl = MUX_s_1_2_2((nor_1273_nl), (nor_1274_nl), acc_2_tmp_7_1[3]);
  assign nor_1268_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[2]))))
      | and_tmp_10);
  assign nor_1269_nl = ~(and_2691_cse | and_tmp_10);
  assign mux_239_nl = MUX_s_1_2_2((nor_1268_nl), (nor_1269_nl), acc_2_tmp_7_1[3]);
  assign mux_240_nl = MUX_s_1_2_2((~ (MAC_LOOP_mux_11_tmp[3])), (MAC_LOOP_mux_11_tmp[3]),
      MAC_LOOP_mux_11_tmp[0]);
  assign nor_1262_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5])
      | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[3])))) | and_tmp_12);
  assign nor_1263_nl = ~(and_2667_cse | and_tmp_12);
  assign mux_242_nl = MUX_s_1_2_2((nor_1262_nl), (nor_1263_nl), acc_2_tmp_7_1[1]);
  assign nor_1260_nl = ~(((~ (acc_2_tmp_7_1[3])) & (acc_2_tmp_7_1[0]) & (acc_2_tmp_7_1[6])
      & (acc_2_tmp_7_1[5]) & (acc_2_tmp_7_1[4]) & (acc_2_tmp_7_1[2])) | and_tmp_13);
  assign nor_1261_nl = ~(and_2667_cse | and_tmp_13);
  assign mux_244_nl = MUX_s_1_2_2((nor_1260_nl), (nor_1261_nl), acc_2_tmp_7_1[1]);
  assign nor_1256_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5])
      | (acc_2_tmp_7_1[6]) | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[3])))) |
      and_tmp_14);
  assign nor_1257_nl = ~(and_2667_cse | and_tmp_14);
  assign mux_246_nl = MUX_s_1_2_2((nor_1256_nl), (nor_1257_nl), acc_2_tmp_7_1[1]);
  assign nor_1253_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[6]))
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[2]))))
      | and_tmp_15);
  assign nor_1254_nl = ~(and_2667_cse | and_tmp_15);
  assign mux_248_nl = MUX_s_1_2_2((nor_1253_nl), (nor_1254_nl), acc_2_tmp_7_1[1]);
  assign nor_1248_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[3])))) |
      and_tmp_16);
  assign nor_1249_nl = ~(and_2671_cse | and_tmp_16);
  assign mux_250_nl = MUX_s_1_2_2((nor_1248_nl), (nor_1249_nl), acc_2_tmp_7_1[2]);
  assign nor_1245_nl = ~(((~ (acc_2_tmp_7_1[3])) & (acc_2_tmp_7_1[0]) & (acc_2_tmp_7_1[6])
      & (acc_2_tmp_7_1[5]) & (acc_2_tmp_7_1[4]) & (acc_2_tmp_7_1[1])) | and_tmp_17);
  assign nor_1246_nl = ~(and_2671_cse | and_tmp_17);
  assign mux_252_nl = MUX_s_1_2_2((nor_1245_nl), (nor_1246_nl), acc_2_tmp_7_1[2]);
  assign nor_1241_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[3]))))
      | and_tmp_18);
  assign nor_1242_nl = ~(and_2671_cse | and_tmp_18);
  assign mux_254_nl = MUX_s_1_2_2((nor_1241_nl), (nor_1242_nl), acc_2_tmp_7_1[2]);
  assign nor_1237_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[6]))
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_19);
  assign nor_1238_nl = ~(and_2671_cse | and_tmp_19);
  assign mux_256_nl = MUX_s_1_2_2((nor_1237_nl), (nor_1238_nl), acc_2_tmp_7_1[2]);
  assign nor_1232_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[3])))) |
      and_tmp_20);
  assign nor_1233_nl = ~(and_2667_cse | and_tmp_20);
  assign mux_258_nl = MUX_s_1_2_2((nor_1232_nl), (nor_1233_nl), acc_2_tmp_7_1[1]);
  assign nor_1228_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[6])) | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[4]))))
      | and_tmp_21);
  assign nor_1229_nl = ~(and_2667_cse | and_tmp_21);
  assign mux_260_nl = MUX_s_1_2_2((nor_1228_nl), (nor_1229_nl), acc_2_tmp_7_1[1]);
  assign nor_1224_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[3]))))
      | and_tmp_22);
  assign nor_1225_nl = ~(and_2667_cse | and_tmp_22);
  assign mux_262_nl = MUX_s_1_2_2((nor_1224_nl), (nor_1225_nl), acc_2_tmp_7_1[1]);
  assign nor_1220_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[6])) | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[4]))))
      | and_tmp_23);
  assign nor_1221_nl = ~(and_2667_cse | and_tmp_23);
  assign mux_264_nl = MUX_s_1_2_2((nor_1220_nl), (nor_1221_nl), acc_2_tmp_7_1[1]);
  assign nor_1215_nl = ~((~((acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_24);
  assign nor_1216_nl = ~(and_2736_cse | and_tmp_24);
  assign mux_266_nl = MUX_s_1_2_2((nor_1215_nl), (nor_1216_nl), acc_2_tmp_7_1[4]);
  assign nor_1210_nl = ~((~((acc_2_tmp_7_1[5:0]!=6'b001111))) | and_tmp_25);
  assign nor_1211_nl = ~(and_2741_cse | and_tmp_25);
  assign mux_268_nl = MUX_s_1_2_2((nor_1210_nl), (nor_1211_nl), acc_2_tmp_7_1[6]);
  assign or_1206_nl = (acc_2_tmp_7_1[4]) | (~ (acc_2_tmp_7_1[0])) | and_tmp_26;
  assign mux_270_nl = MUX_s_1_2_2(and_tmp_26, (or_1206_nl), and_2736_cse);
  assign nor_1205_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[5])
      | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[4])))) | and_tmp_27);
  assign nor_1206_nl = ~(and_2667_cse | and_tmp_27);
  assign mux_272_nl = MUX_s_1_2_2((nor_1205_nl), (nor_1206_nl), acc_2_tmp_7_1[1]);
  assign nor_1203_nl = ~(((~ (acc_2_tmp_7_1[4])) & (acc_2_tmp_7_1[0]) & (acc_2_tmp_7_1[6])
      & (acc_2_tmp_7_1[5]) & (acc_2_tmp_7_1[3]) & (acc_2_tmp_7_1[2])) | and_tmp_28);
  assign nor_1204_nl = ~(and_2667_cse | and_tmp_28);
  assign mux_274_nl = MUX_s_1_2_2((nor_1203_nl), (nor_1204_nl), acc_2_tmp_7_1[1]);
  assign nor_1199_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[5])
      | (acc_2_tmp_7_1[6]) | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[4])))) |
      and_tmp_29);
  assign nor_1200_nl = ~(and_2667_cse | and_tmp_29);
  assign mux_276_nl = MUX_s_1_2_2((nor_1199_nl), (nor_1200_nl), acc_2_tmp_7_1[1]);
  assign nor_1196_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[6]))
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[2]))))
      | and_tmp_30);
  assign nor_1197_nl = ~(and_2667_cse | and_tmp_30);
  assign mux_278_nl = MUX_s_1_2_2((nor_1196_nl), (nor_1197_nl), acc_2_tmp_7_1[1]);
  assign nor_1191_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[4])))) |
      and_tmp_31);
  assign nor_1192_nl = ~(and_2671_cse | and_tmp_31);
  assign mux_280_nl = MUX_s_1_2_2((nor_1191_nl), (nor_1192_nl), acc_2_tmp_7_1[2]);
  assign nor_1189_nl = ~(((~ (acc_2_tmp_7_1[2])) & (acc_2_tmp_7_1[0]) & (acc_2_tmp_7_1[6])
      & (acc_2_tmp_7_1[5]) & (acc_2_tmp_7_1[3]) & (acc_2_tmp_7_1[1])) | and_tmp_32);
  assign nor_1190_nl = ~(and_2736_cse | and_tmp_32);
  assign mux_282_nl = MUX_s_1_2_2((nor_1189_nl), (nor_1190_nl), acc_2_tmp_7_1[4]);
  assign nor_1185_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[4]))))
      | and_tmp_33);
  assign nor_1186_nl = ~(and_2671_cse | and_tmp_33);
  assign mux_284_nl = MUX_s_1_2_2((nor_1185_nl), (nor_1186_nl), acc_2_tmp_7_1[2]);
  assign nor_1182_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[6]))
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_34);
  assign nor_1183_nl = ~(and_2671_cse | and_tmp_34);
  assign mux_286_nl = MUX_s_1_2_2((nor_1182_nl), (nor_1183_nl), acc_2_tmp_7_1[2]);
  assign nor_1178_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[2])))) |
      and_tmp_35);
  assign nor_1179_nl = ~(and_2667_cse | and_tmp_35);
  assign mux_288_nl = MUX_s_1_2_2((nor_1178_nl), (nor_1179_nl), acc_2_tmp_7_1[1]);
  assign nor_1175_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[4]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[6]))))
      | and_tmp_36);
  assign nor_1176_nl = ~(and_2667_cse | and_tmp_36);
  assign mux_290_nl = MUX_s_1_2_2((nor_1175_nl), (nor_1176_nl), acc_2_tmp_7_1[1]);
  assign nor_1172_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[2]))))
      | and_tmp_37);
  assign nor_1173_nl = ~(and_2667_cse | and_tmp_37);
  assign mux_292_nl = MUX_s_1_2_2((nor_1172_nl), (nor_1173_nl), acc_2_tmp_7_1[1]);
  assign nor_1169_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[6]))))
      | and_tmp_38);
  assign nor_1170_nl = ~(and_2667_cse | and_tmp_38);
  assign mux_294_nl = MUX_s_1_2_2((nor_1169_nl), (nor_1170_nl), acc_2_tmp_7_1[1]);
  assign nor_1165_nl = ~((~((acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[4]))))
      | and_tmp_39);
  assign nor_1166_nl = ~(and_2691_cse | and_tmp_39);
  assign mux_296_nl = MUX_s_1_2_2((nor_1165_nl), (nor_1166_nl), acc_2_tmp_7_1[3]);
  assign nor_1163_nl = ~(((~ (acc_2_tmp_7_1[4])) & (acc_2_tmp_7_1[0]) & (acc_2_tmp_7_1[6])
      & (acc_2_tmp_7_1[5]) & (acc_2_tmp_7_1[2]) & (acc_2_tmp_7_1[1])) | and_tmp_40);
  assign nor_1164_nl = ~(and_2691_cse | and_tmp_40);
  assign mux_298_nl = MUX_s_1_2_2((nor_1163_nl), (nor_1164_nl), acc_2_tmp_7_1[3]);
  assign nor_1160_nl = ~((~((acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[4]))))
      | and_tmp_41);
  assign nor_1161_nl = ~(and_2691_cse | and_tmp_41);
  assign mux_300_nl = MUX_s_1_2_2((nor_1160_nl), (nor_1161_nl), acc_2_tmp_7_1[3]);
  assign nor_1157_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[6]))
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_42);
  assign nor_1158_nl = ~(and_2691_cse | and_tmp_42);
  assign mux_302_nl = MUX_s_1_2_2((nor_1157_nl), (nor_1158_nl), acc_2_tmp_7_1[3]);
  assign nor_1153_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[4])))) |
      and_tmp_43);
  assign nor_1154_nl = ~(and_2667_cse | and_tmp_43);
  assign mux_304_nl = MUX_s_1_2_2((nor_1153_nl), (nor_1154_nl), acc_2_tmp_7_1[1]);
  assign nor_1150_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[6]))))
      | and_tmp_44);
  assign nor_1151_nl = ~(and_2667_cse | and_tmp_44);
  assign mux_306_nl = MUX_s_1_2_2((nor_1150_nl), (nor_1151_nl), acc_2_tmp_7_1[1]);
  assign nor_1147_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[4]))))
      | and_tmp_45);
  assign nor_1148_nl = ~(and_2667_cse | and_tmp_45);
  assign mux_308_nl = MUX_s_1_2_2((nor_1147_nl), (nor_1148_nl), acc_2_tmp_7_1[1]);
  assign nor_1144_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[6]))))
      | and_tmp_46);
  assign nor_1145_nl = ~(and_2667_cse | and_tmp_46);
  assign mux_310_nl = MUX_s_1_2_2((nor_1144_nl), (nor_1145_nl), acc_2_tmp_7_1[1]);
  assign nor_1140_nl = ~((~((acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[4]))))
      | and_tmp_47);
  assign nor_1141_nl = ~(and_2671_cse | and_tmp_47);
  assign mux_312_nl = MUX_s_1_2_2((nor_1140_nl), (nor_1141_nl), acc_2_tmp_7_1[2]);
  assign nor_1136_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[2]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[6])) | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_48);
  assign nor_1137_nl = ~(and_2736_cse | and_tmp_48);
  assign mux_314_nl = MUX_s_1_2_2((nor_1136_nl), (nor_1137_nl), acc_2_tmp_7_1[4]);
  assign nor_1133_nl = ~((~((acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[4]))))
      | and_tmp_49);
  assign nor_1134_nl = ~(and_2671_cse | and_tmp_49);
  assign mux_316_nl = MUX_s_1_2_2((nor_1133_nl), (nor_1134_nl), acc_2_tmp_7_1[2]);
  assign nor_1129_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[6])) | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_50);
  assign nor_1130_nl = ~(and_2671_cse | and_tmp_50);
  assign mux_318_nl = MUX_s_1_2_2((nor_1129_nl), (nor_1130_nl), acc_2_tmp_7_1[2]);
  assign nor_1125_nl = ~((~((acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[2]))))
      | and_tmp_51);
  assign nor_1126_nl = ~(and_2667_cse | and_tmp_51);
  assign mux_320_nl = MUX_s_1_2_2((nor_1125_nl), (nor_1126_nl), acc_2_tmp_7_1[1]);
  assign nor_1121_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[6]))))
      | and_tmp_52);
  assign nor_1122_nl = ~(and_2667_cse | and_tmp_52);
  assign mux_322_nl = MUX_s_1_2_2((nor_1121_nl), (nor_1122_nl), acc_2_tmp_7_1[1]);
  assign nor_1118_nl = ~((~((acc_2_tmp_7_1[5:0]!=6'b011101))) | and_tmp_53);
  assign nor_1119_nl = ~(and_2741_cse | and_tmp_53);
  assign mux_324_nl = MUX_s_1_2_2((nor_1118_nl), (nor_1119_nl), acc_2_tmp_7_1[6]);
  assign nor_1114_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[6])))) |
      and_tmp_54);
  assign nor_1115_nl = ~(and_2667_cse | and_tmp_54);
  assign mux_326_nl = MUX_s_1_2_2((nor_1114_nl), (nor_1115_nl), acc_2_tmp_7_1[1]);
  assign nor_1110_nl = ~((~((acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[4]))
      | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_55);
  assign nor_1111_nl = ~(and_2829_cse | and_tmp_55);
  assign mux_328_nl = MUX_s_1_2_2((nor_1110_nl), (nor_1111_nl), acc_2_tmp_7_1[5]);
  assign nor_1107_nl = ~(((~ (acc_2_tmp_7_1[6])) & (acc_2_tmp_7_1[0]) & (acc_2_tmp_7_1[4])
      & (acc_2_tmp_7_1[3]) & (acc_2_tmp_7_1[2]) & (acc_2_tmp_7_1[1])) | and_tmp_56);
  assign nor_1108_nl = ~(and_2829_cse | and_tmp_56);
  assign mux_330_nl = MUX_s_1_2_2((nor_1107_nl), (nor_1108_nl), acc_2_tmp_7_1[5]);
  assign or_1205_nl = (acc_2_tmp_7_1[5]) | (~ (acc_2_tmp_7_1[0])) | and_tmp_57;
  assign mux_332_nl = MUX_s_1_2_2(and_tmp_57, (or_1205_nl), and_2829_cse);
  assign nor_1101_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4])
      | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[5])))) | and_tmp_58);
  assign nor_1102_nl = ~(and_2667_cse | and_tmp_58);
  assign mux_334_nl = MUX_s_1_2_2((nor_1101_nl), (nor_1102_nl), acc_2_tmp_7_1[1]);
  assign nor_1099_nl = ~(((~ (acc_2_tmp_7_1[5])) & (acc_2_tmp_7_1[0]) & (acc_2_tmp_7_1[6])
      & (acc_2_tmp_7_1[4]) & (acc_2_tmp_7_1[3]) & (acc_2_tmp_7_1[2])) | and_tmp_59);
  assign nor_1100_nl = ~(and_2667_cse | and_tmp_59);
  assign mux_336_nl = MUX_s_1_2_2((nor_1099_nl), (nor_1100_nl), acc_2_tmp_7_1[1]);
  assign nor_1094_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4])
      | (acc_2_tmp_7_1[6]) | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[5])))) |
      and_tmp_60);
  assign nor_1095_nl = ~(and_2667_cse | and_tmp_60);
  assign mux_338_nl = MUX_s_1_2_2((nor_1094_nl), (nor_1095_nl), acc_2_tmp_7_1[1]);
  assign nor_1090_nl = ~((~((acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[6]))
      | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[2]))))
      | and_tmp_61);
  assign nor_1091_nl = ~(and_2667_cse | and_tmp_61);
  assign mux_340_nl = MUX_s_1_2_2((nor_1090_nl), (nor_1091_nl), acc_2_tmp_7_1[1]);
  assign nor_1085_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[6])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[5])))) |
      and_tmp_62);
  assign nor_1086_nl = ~(and_2671_cse | and_tmp_62);
  assign mux_342_nl = MUX_s_1_2_2((nor_1085_nl), (nor_1086_nl), acc_2_tmp_7_1[2]);
  assign nor_1083_nl = ~(((~ (acc_2_tmp_7_1[5])) & (acc_2_tmp_7_1[0]) & (acc_2_tmp_7_1[6])
      & (acc_2_tmp_7_1[1]) & (acc_2_tmp_7_1[3]) & (acc_2_tmp_7_1[4])) | and_tmp_63);
  assign nor_1084_nl = ~(and_2671_cse | and_tmp_63);
  assign mux_344_nl = MUX_s_1_2_2((nor_1083_nl), (nor_1084_nl), acc_2_tmp_7_1[2]);
  assign nor_1078_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[6])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[5]))))
      | and_tmp_64);
  assign nor_1079_nl = ~(and_2671_cse | and_tmp_64);
  assign mux_346_nl = MUX_s_1_2_2((nor_1078_nl), (nor_1079_nl), acc_2_tmp_7_1[2]);
  assign nor_1074_nl = ~((~((acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[6]))
      | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[4]))))
      | and_tmp_65);
  assign nor_1075_nl = ~(and_2671_cse | and_tmp_65);
  assign mux_348_nl = MUX_s_1_2_2((nor_1074_nl), (nor_1075_nl), acc_2_tmp_7_1[2]);
  assign nor_1070_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[6])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[5])))) |
      and_tmp_66);
  assign nor_1071_nl = ~(and_2667_cse | and_tmp_66);
  assign mux_350_nl = MUX_s_1_2_2((nor_1070_nl), (nor_1071_nl), acc_2_tmp_7_1[1]);
  assign nor_1067_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[1]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[6]))))
      | and_tmp_67);
  assign nor_1068_nl = ~(and_2829_cse | and_tmp_67);
  assign mux_352_nl = MUX_s_1_2_2((nor_1067_nl), (nor_1068_nl), acc_2_tmp_7_1[5]);
  assign nor_1063_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[6])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[5]))))
      | and_tmp_68);
  assign nor_1064_nl = ~(and_2667_cse | and_tmp_68);
  assign mux_354_nl = MUX_s_1_2_2((nor_1063_nl), (nor_1064_nl), acc_2_tmp_7_1[1]);
  assign nor_1059_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[6]))))
      | and_tmp_69);
  assign nor_1060_nl = ~(and_2667_cse | and_tmp_69);
  assign mux_356_nl = MUX_s_1_2_2((nor_1059_nl), (nor_1060_nl), acc_2_tmp_7_1[1]);
  assign nor_1055_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_70);
  assign nor_1056_nl = ~(and_2691_cse | and_tmp_70);
  assign mux_358_nl = MUX_s_1_2_2((nor_1055_nl), (nor_1056_nl), acc_2_tmp_7_1[3]);
  assign nor_1053_nl = ~(((~ (acc_2_tmp_7_1[5])) & (acc_2_tmp_7_1[0]) & (acc_2_tmp_7_1[6])
      & (acc_2_tmp_7_1[1]) & (acc_2_tmp_7_1[2]) & (acc_2_tmp_7_1[4])) | and_tmp_71);
  assign nor_1054_nl = ~(and_2691_cse | and_tmp_71);
  assign mux_360_nl = MUX_s_1_2_2((nor_1053_nl), (nor_1054_nl), acc_2_tmp_7_1[3]);
  assign nor_1049_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[6]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_72);
  assign nor_1050_nl = ~(and_2691_cse | and_tmp_72);
  assign mux_362_nl = MUX_s_1_2_2((nor_1049_nl), (nor_1050_nl), acc_2_tmp_7_1[3]);
  assign nor_1045_nl = ~((~((acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[6]))
      | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[4]))))
      | and_tmp_73);
  assign nor_1046_nl = ~(and_2691_cse | and_tmp_73);
  assign mux_364_nl = MUX_s_1_2_2((nor_1045_nl), (nor_1046_nl), acc_2_tmp_7_1[3]);
  assign nor_1041_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[6])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[5])))) |
      and_tmp_74);
  assign nor_1042_nl = ~(and_2667_cse | and_tmp_74);
  assign mux_366_nl = MUX_s_1_2_2((nor_1041_nl), (nor_1042_nl), acc_2_tmp_7_1[1]);
  assign nor_1038_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[1]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[6]))))
      | and_tmp_75);
  assign nor_1039_nl = ~(and_2829_cse | and_tmp_75);
  assign mux_368_nl = MUX_s_1_2_2((nor_1038_nl), (nor_1039_nl), acc_2_tmp_7_1[5]);
  assign nor_1034_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[6])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[5]))))
      | and_tmp_76);
  assign nor_1035_nl = ~(and_2667_cse | and_tmp_76);
  assign mux_370_nl = MUX_s_1_2_2((nor_1034_nl), (nor_1035_nl), acc_2_tmp_7_1[1]);
  assign nor_1030_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[6]))))
      | and_tmp_77);
  assign nor_1031_nl = ~(and_2667_cse | and_tmp_77);
  assign mux_372_nl = MUX_s_1_2_2((nor_1030_nl), (nor_1031_nl), acc_2_tmp_7_1[1]);
  assign nor_1026_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_78);
  assign nor_1027_nl = ~(and_2671_cse | and_tmp_78);
  assign mux_374_nl = MUX_s_1_2_2((nor_1026_nl), (nor_1027_nl), acc_2_tmp_7_1[2]);
  assign nor_1022_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[2]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[6])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_79);
  assign nor_1023_nl = ~(and_2829_cse | and_tmp_79);
  assign mux_376_nl = MUX_s_1_2_2((nor_1022_nl), (nor_1023_nl), acc_2_tmp_7_1[5]);
  assign nor_1018_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[6]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_80);
  assign nor_1019_nl = ~(and_2671_cse | and_tmp_80);
  assign mux_378_nl = MUX_s_1_2_2((nor_1018_nl), (nor_1019_nl), acc_2_tmp_7_1[2]);
  assign nor_1013_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[6])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_81);
  assign nor_1014_nl = ~(and_2671_cse | and_tmp_81);
  assign mux_380_nl = MUX_s_1_2_2((nor_1013_nl), (nor_1014_nl), acc_2_tmp_7_1[2]);
  assign nor_1009_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[2]))))
      | and_tmp_82);
  assign nor_1010_nl = ~(and_2667_cse | and_tmp_82);
  assign mux_382_nl = MUX_s_1_2_2((nor_1009_nl), (nor_1010_nl), acc_2_tmp_7_1[1]);
  assign nor_1005_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[5])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[6])) | (~ (acc_2_tmp_7_1[4]))))
      | and_tmp_83);
  assign nor_1006_nl = ~(and_2667_cse | and_tmp_83);
  assign mux_384_nl = MUX_s_1_2_2((nor_1005_nl), (nor_1006_nl), acc_2_tmp_7_1[1]);
  assign nor_1001_nl = ~((~((acc_2_tmp_7_1[5:0]!=6'b101101))) | and_tmp_84);
  assign nor_1002_nl = ~(and_2741_cse | and_tmp_84);
  assign mux_386_nl = MUX_s_1_2_2((nor_1001_nl), (nor_1002_nl), acc_2_tmp_7_1[6]);
  assign nor_996_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[5])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[6])) | (~ (acc_2_tmp_7_1[4])))) |
      and_tmp_85);
  assign nor_997_nl = ~(and_2667_cse | and_tmp_85);
  assign mux_388_nl = MUX_s_1_2_2((nor_996_nl), (nor_997_nl), acc_2_tmp_7_1[1]);
  assign nor_992_nl = ~((~((acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[5]))
      | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_86);
  assign nor_993_nl = ~(and_2736_cse | and_tmp_86);
  assign mux_390_nl = MUX_s_1_2_2((nor_992_nl), (nor_993_nl), acc_2_tmp_7_1[4]);
  assign nor_990_nl = ~(((~ (acc_2_tmp_7_1[5])) & (acc_2_tmp_7_1[0]) & (acc_2_tmp_7_1[6])
      & (acc_2_tmp_7_1[3]) & (acc_2_tmp_7_1[2]) & (acc_2_tmp_7_1[1])) | and_tmp_87);
  assign nor_991_nl = ~(and_2736_cse | and_tmp_87);
  assign mux_392_nl = MUX_s_1_2_2((nor_990_nl), (nor_991_nl), acc_2_tmp_7_1[4]);
  assign nor_987_nl = ~(((acc_2_tmp_7_1[5:0]==6'b101111)) | and_tmp_88);
  assign nor_988_nl = ~(and_2741_cse | and_tmp_88);
  assign mux_394_nl = MUX_s_1_2_2((nor_987_nl), (nor_988_nl), acc_2_tmp_7_1[6]);
  assign nor_983_nl = ~((~((acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[6]))
      | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_89);
  assign nor_984_nl = ~(and_2736_cse | and_tmp_89);
  assign mux_396_nl = MUX_s_1_2_2((nor_983_nl), (nor_984_nl), acc_2_tmp_7_1[4]);
  assign nor_979_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[6])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[5])))) |
      and_tmp_90);
  assign nor_980_nl = ~(and_2667_cse | and_tmp_90);
  assign mux_398_nl = MUX_s_1_2_2((nor_979_nl), (nor_980_nl), acc_2_tmp_7_1[1]);
  assign nor_976_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[1]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[6]))))
      | and_tmp_91);
  assign nor_977_nl = ~(and_2829_cse | and_tmp_91);
  assign mux_400_nl = MUX_s_1_2_2((nor_976_nl), (nor_977_nl), acc_2_tmp_7_1[5]);
  assign nor_972_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[6])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[5]))))
      | and_tmp_92);
  assign nor_973_nl = ~(and_2667_cse | and_tmp_92);
  assign mux_402_nl = MUX_s_1_2_2((nor_972_nl), (nor_973_nl), acc_2_tmp_7_1[1]);
  assign nor_968_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[6]))))
      | and_tmp_93);
  assign nor_969_nl = ~(and_2667_cse | and_tmp_93);
  assign mux_404_nl = MUX_s_1_2_2((nor_968_nl), (nor_969_nl), acc_2_tmp_7_1[1]);
  assign nor_964_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_94);
  assign nor_965_nl = ~(and_2671_cse | and_tmp_94);
  assign mux_406_nl = MUX_s_1_2_2((nor_964_nl), (nor_965_nl), acc_2_tmp_7_1[2]);
  assign nor_961_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[2]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[6])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_95);
  assign nor_962_nl = ~(and_2829_cse | and_tmp_95);
  assign mux_408_nl = MUX_s_1_2_2((nor_961_nl), (nor_962_nl), acc_2_tmp_7_1[5]);
  assign nor_957_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[6]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_96);
  assign nor_958_nl = ~(and_2671_cse | and_tmp_96);
  assign mux_410_nl = MUX_s_1_2_2((nor_957_nl), (nor_958_nl), acc_2_tmp_7_1[2]);
  assign nor_953_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[6])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_97);
  assign nor_954_nl = ~(and_2671_cse | and_tmp_97);
  assign mux_412_nl = MUX_s_1_2_2((nor_953_nl), (nor_954_nl), acc_2_tmp_7_1[2]);
  assign nor_950_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[2]))))
      | and_tmp_98);
  assign nor_951_nl = ~(and_2667_cse | and_tmp_98);
  assign mux_414_nl = MUX_s_1_2_2((nor_950_nl), (nor_951_nl), acc_2_tmp_7_1[1]);
  assign nor_947_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[6]))))
      | and_tmp_99);
  assign nor_948_nl = ~(and_2667_cse | and_tmp_99);
  assign mux_416_nl = MUX_s_1_2_2((nor_947_nl), (nor_948_nl), acc_2_tmp_7_1[1]);
  assign nor_944_nl = ~((~((acc_2_tmp_7_1[5:0]!=6'b110101))) | and_tmp_100);
  assign nor_945_nl = ~(and_2741_cse | and_tmp_100);
  assign mux_418_nl = MUX_s_1_2_2((nor_944_nl), (nor_945_nl), acc_2_tmp_7_1[6]);
  assign nor_940_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[6])))) |
      and_tmp_101);
  assign nor_941_nl = ~(and_2667_cse | and_tmp_101);
  assign mux_420_nl = MUX_s_1_2_2((nor_940_nl), (nor_941_nl), acc_2_tmp_7_1[1]);
  assign nor_937_nl = ~((~((acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[5]))
      | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[4]))))
      | and_tmp_102);
  assign nor_938_nl = ~(and_2691_cse | and_tmp_102);
  assign mux_422_nl = MUX_s_1_2_2((nor_937_nl), (nor_938_nl), acc_2_tmp_7_1[3]);
  assign nor_934_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[3]) | (~ (acc_2_tmp_7_1[0]))
      | (~ (acc_2_tmp_7_1[6])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_103);
  assign nor_935_nl = ~(and_2829_cse | and_tmp_103);
  assign mux_424_nl = MUX_s_1_2_2((nor_934_nl), (nor_935_nl), acc_2_tmp_7_1[5]);
  assign nor_932_nl = ~(((~ (acc_2_tmp_7_1[6])) & (acc_2_tmp_7_1[0]) & (acc_2_tmp_7_1[5])
      & (acc_2_tmp_7_1[1]) & (acc_2_tmp_7_1[2]) & (acc_2_tmp_7_1[4])) | and_tmp_104);
  assign nor_933_nl = ~(and_2691_cse | and_tmp_104);
  assign mux_426_nl = MUX_s_1_2_2((nor_932_nl), (nor_933_nl), acc_2_tmp_7_1[3]);
  assign nor_928_nl = ~((~((acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[6])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_105);
  assign nor_929_nl = ~(and_2691_cse | and_tmp_105);
  assign mux_428_nl = MUX_s_1_2_2((nor_928_nl), (nor_929_nl), acc_2_tmp_7_1[3]);
  assign nor_925_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0])
      | (~ (acc_2_tmp_7_1[5])) | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[3]))))
      | and_tmp_106);
  assign nor_926_nl = ~(and_2667_cse | and_tmp_106);
  assign mux_430_nl = MUX_s_1_2_2((nor_925_nl), (nor_926_nl), acc_2_tmp_7_1[1]);
  assign nor_922_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[6]))))
      | and_tmp_107);
  assign nor_923_nl = ~(and_2667_cse | and_tmp_107);
  assign mux_432_nl = MUX_s_1_2_2((nor_922_nl), (nor_923_nl), acc_2_tmp_7_1[1]);
  assign nor_919_nl = ~((~((acc_2_tmp_7_1[5:0]!=6'b111001))) | and_tmp_108);
  assign nor_920_nl = ~(and_2741_cse | and_tmp_108);
  assign mux_434_nl = MUX_s_1_2_2((nor_919_nl), (nor_920_nl), acc_2_tmp_7_1[6]);
  assign nor_915_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[2])) | (~ (acc_2_tmp_7_1[6])))) |
      and_tmp_109);
  assign nor_916_nl = ~(and_2667_cse | and_tmp_109);
  assign mux_436_nl = MUX_s_1_2_2((nor_915_nl), (nor_916_nl), acc_2_tmp_7_1[1]);
  assign nor_912_nl = ~((~((acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[5]))
      | (~ (acc_2_tmp_7_1[1])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[4]))))
      | and_tmp_110);
  assign nor_913_nl = ~(and_2671_cse | and_tmp_110);
  assign mux_438_nl = MUX_s_1_2_2((nor_912_nl), (nor_913_nl), acc_2_tmp_7_1[2]);
  assign nor_908_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5])
      | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[6])) | (~ (acc_2_tmp_7_1[1]))))
      | and_tmp_111);
  assign nor_909_nl = ~(and_2671_cse | and_tmp_111);
  assign mux_440_nl = MUX_s_1_2_2((nor_908_nl), (nor_909_nl), acc_2_tmp_7_1[2]);
  assign nor_906_nl = ~(((~ (acc_2_tmp_7_1[6])) & (acc_2_tmp_7_1[0]) & (acc_2_tmp_7_1[5])
      & (acc_2_tmp_7_1[1]) & (acc_2_tmp_7_1[3]) & (acc_2_tmp_7_1[4])) | and_tmp_112);
  assign nor_907_nl = ~(and_2671_cse | and_tmp_112);
  assign mux_442_nl = MUX_s_1_2_2((nor_906_nl), (nor_907_nl), acc_2_tmp_7_1[2]);
  assign nor_901_nl = ~((~((acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4]) | (acc_2_tmp_7_1[5])
      | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[6])) | (~ (acc_2_tmp_7_1[1])))) |
      and_tmp_113);
  assign nor_902_nl = ~(and_2671_cse | and_tmp_113);
  assign mux_444_nl = MUX_s_1_2_2((nor_901_nl), (nor_902_nl), acc_2_tmp_7_1[2]);
  assign nor_898_nl = ~((~((acc_2_tmp_7_1[6]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[5]))
      | (~ (acc_2_tmp_7_1[4])) | (~ (acc_2_tmp_7_1[3])) | (~ (acc_2_tmp_7_1[2]))))
      | and_tmp_114);
  assign nor_899_nl = ~(and_2667_cse | and_tmp_114);
  assign mux_446_nl = MUX_s_1_2_2((nor_898_nl), (nor_899_nl), acc_2_tmp_7_1[1]);
  assign nor_894_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4])
      | (acc_2_tmp_7_1[5]) | (~ (acc_2_tmp_7_1[0])) | (~ (acc_2_tmp_7_1[6])))) |
      and_tmp_115);
  assign nor_895_nl = ~(and_2667_cse | and_tmp_115);
  assign mux_448_nl = MUX_s_1_2_2((nor_894_nl), (nor_895_nl), acc_2_tmp_7_1[1]);
  assign nor_892_nl = ~(((acc_2_tmp_7_1[5:0]==6'b111101)) | and_tmp_116);
  assign nor_893_nl = ~(and_2741_cse | and_tmp_116);
  assign mux_450_nl = MUX_s_1_2_2((nor_892_nl), (nor_893_nl), acc_2_tmp_7_1[6]);
  assign nor_887_nl = ~((~((acc_2_tmp_7_1[2]) | (acc_2_tmp_7_1[3]) | (acc_2_tmp_7_1[4])
      | (acc_2_tmp_7_1[5]) | (acc_2_tmp_7_1[0]) | (~ (acc_2_tmp_7_1[6])))) | and_tmp_117);
  assign nor_888_nl = ~(and_2667_cse | and_tmp_117);
  assign mux_452_nl = MUX_s_1_2_2((nor_887_nl), (nor_888_nl), acc_2_tmp_7_1[1]);
  assign or_1204_nl = (acc_2_tmp_7_1[6]) | (~ (acc_2_tmp_7_1[0])) | and_tmp_118;
  assign mux_454_nl = MUX_s_1_2_2(and_tmp_118, (or_1204_nl), and_2741_cse);
  assign SHIFT_LOOP_n_or_nl = (z_out_1_7 & (fsm_output[1])) | (fsm_output[2]);
  assign SHIFT_LOOP_n_SHIFT_LOOP_n_mux_nl = MUX_v_7_2_2(7'b1111110, acc_2_tmp_7_1,
      SHIFT_LOOP_n_or_nl);
  assign MAC_LOOP_n_nor_nl = ~((fsm_output[4:3]!=2'b00) | ((~ z_out_1_7) & (fsm_output[1])));
  assign SHIFT_LOOP_mux_129_nl = MUX_v_7_2_2((~ acc_2_tmp_7_1), acc_2_tmp_7_1, fsm_output[2]);
  assign nl_SHIFT_LOOP_acc_nl = ({1'b1 , (SHIFT_LOOP_mux_129_nl)}) + 8'b00000001;
  assign SHIFT_LOOP_acc_nl = nl_SHIFT_LOOP_acc_nl[7:0];
  assign z_out_1_7 = readslicef_8_1_7((SHIFT_LOOP_acc_nl));
  assign MAC_LOOP_mux_7_nl = MUX_v_19_2_2((sum_sva[18:0]), (signext_19_14(sum_sva[19:6])),
      fsm_output[3]);
  assign MAC_LOOP_mux_9_nl = MUX_v_10_127_2((b_rsci_idat[9:0]), (b_rsci_idat[19:10]),
      (b_rsci_idat[29:20]), (b_rsci_idat[39:30]), (b_rsci_idat[49:40]), (b_rsci_idat[59:50]),
      (b_rsci_idat[69:60]), (b_rsci_idat[79:70]), (b_rsci_idat[89:80]), (b_rsci_idat[99:90]),
      (b_rsci_idat[109:100]), (b_rsci_idat[119:110]), (b_rsci_idat[129:120]), (b_rsci_idat[139:130]),
      (b_rsci_idat[149:140]), (b_rsci_idat[159:150]), (b_rsci_idat[169:160]), (b_rsci_idat[179:170]),
      (b_rsci_idat[189:180]), (b_rsci_idat[199:190]), (b_rsci_idat[209:200]), (b_rsci_idat[219:210]),
      (b_rsci_idat[229:220]), (b_rsci_idat[239:230]), (b_rsci_idat[249:240]), (b_rsci_idat[259:250]),
      (b_rsci_idat[269:260]), (b_rsci_idat[279:270]), (b_rsci_idat[289:280]), (b_rsci_idat[299:290]),
      (b_rsci_idat[309:300]), (b_rsci_idat[319:310]), (b_rsci_idat[329:320]), (b_rsci_idat[339:330]),
      (b_rsci_idat[349:340]), (b_rsci_idat[359:350]), (b_rsci_idat[369:360]), (b_rsci_idat[379:370]),
      (b_rsci_idat[389:380]), (b_rsci_idat[399:390]), (b_rsci_idat[409:400]), (b_rsci_idat[419:410]),
      (b_rsci_idat[429:420]), (b_rsci_idat[439:430]), (b_rsci_idat[449:440]), (b_rsci_idat[459:450]),
      (b_rsci_idat[469:460]), (b_rsci_idat[479:470]), (b_rsci_idat[489:480]), (b_rsci_idat[499:490]),
      (b_rsci_idat[509:500]), (b_rsci_idat[519:510]), (b_rsci_idat[529:520]), (b_rsci_idat[539:530]),
      (b_rsci_idat[549:540]), (b_rsci_idat[559:550]), (b_rsci_idat[569:560]), (b_rsci_idat[579:570]),
      (b_rsci_idat[589:580]), (b_rsci_idat[599:590]), (b_rsci_idat[609:600]), (b_rsci_idat[619:610]),
      (b_rsci_idat[629:620]), (b_rsci_idat[639:630]), (b_rsci_idat[649:640]), (b_rsci_idat[659:650]),
      (b_rsci_idat[669:660]), (b_rsci_idat[679:670]), (b_rsci_idat[689:680]), (b_rsci_idat[699:690]),
      (b_rsci_idat[709:700]), (b_rsci_idat[719:710]), (b_rsci_idat[729:720]), (b_rsci_idat[739:730]),
      (b_rsci_idat[749:740]), (b_rsci_idat[759:750]), (b_rsci_idat[769:760]), (b_rsci_idat[779:770]),
      (b_rsci_idat[789:780]), (b_rsci_idat[799:790]), (b_rsci_idat[809:800]), (b_rsci_idat[819:810]),
      (b_rsci_idat[829:820]), (b_rsci_idat[839:830]), (b_rsci_idat[849:840]), (b_rsci_idat[859:850]),
      (b_rsci_idat[869:860]), (b_rsci_idat[879:870]), (b_rsci_idat[889:880]), (b_rsci_idat[899:890]),
      (b_rsci_idat[909:900]), (b_rsci_idat[919:910]), (b_rsci_idat[929:920]), (b_rsci_idat[939:930]),
      (b_rsci_idat[949:940]), (b_rsci_idat[959:950]), (b_rsci_idat[969:960]), (b_rsci_idat[979:970]),
      (b_rsci_idat[989:980]), (b_rsci_idat[999:990]), (b_rsci_idat[1009:1000]), (b_rsci_idat[1019:1010]),
      (b_rsci_idat[1029:1020]), (b_rsci_idat[1039:1030]), (b_rsci_idat[1049:1040]),
      (b_rsci_idat[1059:1050]), (b_rsci_idat[1069:1060]), (b_rsci_idat[1079:1070]),
      (b_rsci_idat[1089:1080]), (b_rsci_idat[1099:1090]), (b_rsci_idat[1109:1100]),
      (b_rsci_idat[1119:1110]), (b_rsci_idat[1129:1120]), (b_rsci_idat[1139:1130]),
      (b_rsci_idat[1149:1140]), (b_rsci_idat[1159:1150]), (b_rsci_idat[1169:1160]),
      (b_rsci_idat[1179:1170]), (b_rsci_idat[1189:1180]), (b_rsci_idat[1199:1190]),
      (b_rsci_idat[1209:1200]), (b_rsci_idat[1219:1210]), (b_rsci_idat[1229:1220]),
      (b_rsci_idat[1239:1230]), (b_rsci_idat[1249:1240]), (b_rsci_idat[1259:1250]),
      (b_rsci_idat[1269:1260]), MAC_LOOP_n_6_0_sva);
  assign MAC_LOOP_mul_1_nl = conv_s2u_13_13($signed(z_out) * $signed((MAC_LOOP_mux_9_nl)));
  assign MAC_LOOP_mux_8_nl = MUX_v_13_2_2((MAC_LOOP_mul_1_nl), ({12'b000000000000
      , (sum_sva[5])}), fsm_output[3]);
  assign nl_z_out_2 = ({(sum_sva[19]) , (MAC_LOOP_mux_7_nl)}) + conv_s2u_13_20(MAC_LOOP_mux_8_nl);
  assign z_out_2 = nl_z_out_2[19:0];
  assign nl_acc_2_tmp_7_1 = MAC_LOOP_n_6_0_sva + conv_s2u_2_7({(fsm_output[1]) ,
      1'b1});
  assign acc_2_tmp_7_1 = nl_acc_2_tmp_7_1[6:0];
  assign MAC_LOOP_mux_11_tmp = MUX_v_7_2_2(MAC_LOOP_n_6_0_sva, acc_2_tmp_7_1, fsm_output[1]);
  assign MAC_LOOP_mux_10_nl = MUX_v_3_2_2(i_sample_sva, x_0_sva, fsm_output[1]);
  assign z_out = MUX_v_3_127_2((MAC_LOOP_mux_10_nl), x_1_lpi_2, x_2_lpi_2, x_3_lpi_2,
      x_4_lpi_2, x_5_lpi_2, x_6_lpi_2, x_7_lpi_2, x_8_lpi_2, x_9_lpi_2, x_10_lpi_2,
      x_11_lpi_2, x_12_lpi_2, x_13_lpi_2, x_14_lpi_2, x_15_lpi_2, x_16_lpi_2, x_17_lpi_2,
      x_18_lpi_2, x_19_lpi_2, x_20_lpi_2, x_21_lpi_2, x_22_lpi_2, x_23_lpi_2, x_24_lpi_2,
      x_25_lpi_2, x_26_lpi_2, x_27_lpi_2, x_28_lpi_2, x_29_lpi_2, x_30_lpi_2, x_31_lpi_2,
      x_32_lpi_2, x_33_lpi_2, x_34_lpi_2, x_35_lpi_2, x_36_lpi_2, x_37_lpi_2, x_38_lpi_2,
      x_39_lpi_2, x_40_lpi_2, x_41_lpi_2, x_42_lpi_2, x_43_lpi_2, x_44_lpi_2, x_45_lpi_2,
      x_46_lpi_2, x_47_lpi_2, x_48_lpi_2, x_49_lpi_2, x_50_lpi_2, x_51_lpi_2, x_52_lpi_2,
      x_53_lpi_2, x_54_lpi_2, x_55_lpi_2, x_56_lpi_2, x_57_lpi_2, x_58_lpi_2, x_59_lpi_2,
      x_60_lpi_2, x_61_lpi_2, x_62_lpi_2, x_63_lpi_2, x_64_lpi_2, x_65_lpi_2, x_66_lpi_2,
      x_67_lpi_2, x_68_lpi_2, x_69_lpi_2, x_70_lpi_2, x_71_lpi_2, x_72_lpi_2, x_73_lpi_2,
      x_74_lpi_2, x_75_lpi_2, x_76_lpi_2, x_77_lpi_2, x_78_lpi_2, x_79_lpi_2, x_80_lpi_2,
      x_81_lpi_2, x_82_lpi_2, x_83_lpi_2, x_84_lpi_2, x_85_lpi_2, x_86_lpi_2, x_87_lpi_2,
      x_88_lpi_2, x_89_lpi_2, x_90_lpi_2, x_91_lpi_2, x_92_lpi_2, x_93_lpi_2, x_94_lpi_2,
      x_95_lpi_2, x_96_lpi_2, x_97_lpi_2, x_98_lpi_2, x_99_lpi_2, x_100_lpi_2, x_101_lpi_2,
      x_102_lpi_2, x_103_lpi_2, x_104_lpi_2, x_105_lpi_2, x_106_lpi_2, x_107_lpi_2,
      x_108_lpi_2, x_109_lpi_2, x_110_lpi_2, x_111_lpi_2, x_112_lpi_2, x_113_lpi_2,
      x_114_lpi_2, x_115_lpi_2, x_116_lpi_2, x_117_lpi_2, x_118_lpi_2, x_119_lpi_2,
      x_120_lpi_2, x_121_lpi_2, x_122_lpi_2, x_123_lpi_2, x_124_lpi_2, x_125_lpi_2,
      x_126_lpi_2, MAC_LOOP_mux_11_tmp);

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_127_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input [9:0] input_2;
    input [9:0] input_3;
    input [9:0] input_4;
    input [9:0] input_5;
    input [9:0] input_6;
    input [9:0] input_7;
    input [9:0] input_8;
    input [9:0] input_9;
    input [9:0] input_10;
    input [9:0] input_11;
    input [9:0] input_12;
    input [9:0] input_13;
    input [9:0] input_14;
    input [9:0] input_15;
    input [9:0] input_16;
    input [9:0] input_17;
    input [9:0] input_18;
    input [9:0] input_19;
    input [9:0] input_20;
    input [9:0] input_21;
    input [9:0] input_22;
    input [9:0] input_23;
    input [9:0] input_24;
    input [9:0] input_25;
    input [9:0] input_26;
    input [9:0] input_27;
    input [9:0] input_28;
    input [9:0] input_29;
    input [9:0] input_30;
    input [9:0] input_31;
    input [9:0] input_32;
    input [9:0] input_33;
    input [9:0] input_34;
    input [9:0] input_35;
    input [9:0] input_36;
    input [9:0] input_37;
    input [9:0] input_38;
    input [9:0] input_39;
    input [9:0] input_40;
    input [9:0] input_41;
    input [9:0] input_42;
    input [9:0] input_43;
    input [9:0] input_44;
    input [9:0] input_45;
    input [9:0] input_46;
    input [9:0] input_47;
    input [9:0] input_48;
    input [9:0] input_49;
    input [9:0] input_50;
    input [9:0] input_51;
    input [9:0] input_52;
    input [9:0] input_53;
    input [9:0] input_54;
    input [9:0] input_55;
    input [9:0] input_56;
    input [9:0] input_57;
    input [9:0] input_58;
    input [9:0] input_59;
    input [9:0] input_60;
    input [9:0] input_61;
    input [9:0] input_62;
    input [9:0] input_63;
    input [9:0] input_64;
    input [9:0] input_65;
    input [9:0] input_66;
    input [9:0] input_67;
    input [9:0] input_68;
    input [9:0] input_69;
    input [9:0] input_70;
    input [9:0] input_71;
    input [9:0] input_72;
    input [9:0] input_73;
    input [9:0] input_74;
    input [9:0] input_75;
    input [9:0] input_76;
    input [9:0] input_77;
    input [9:0] input_78;
    input [9:0] input_79;
    input [9:0] input_80;
    input [9:0] input_81;
    input [9:0] input_82;
    input [9:0] input_83;
    input [9:0] input_84;
    input [9:0] input_85;
    input [9:0] input_86;
    input [9:0] input_87;
    input [9:0] input_88;
    input [9:0] input_89;
    input [9:0] input_90;
    input [9:0] input_91;
    input [9:0] input_92;
    input [9:0] input_93;
    input [9:0] input_94;
    input [9:0] input_95;
    input [9:0] input_96;
    input [9:0] input_97;
    input [9:0] input_98;
    input [9:0] input_99;
    input [9:0] input_100;
    input [9:0] input_101;
    input [9:0] input_102;
    input [9:0] input_103;
    input [9:0] input_104;
    input [9:0] input_105;
    input [9:0] input_106;
    input [9:0] input_107;
    input [9:0] input_108;
    input [9:0] input_109;
    input [9:0] input_110;
    input [9:0] input_111;
    input [9:0] input_112;
    input [9:0] input_113;
    input [9:0] input_114;
    input [9:0] input_115;
    input [9:0] input_116;
    input [9:0] input_117;
    input [9:0] input_118;
    input [9:0] input_119;
    input [9:0] input_120;
    input [9:0] input_121;
    input [9:0] input_122;
    input [9:0] input_123;
    input [9:0] input_124;
    input [9:0] input_125;
    input [9:0] input_126;
    input [6:0] sel;
    reg [9:0] result;
  begin
    case (sel)
      7'b0000000 : begin
        result = input_0;
      end
      7'b0000001 : begin
        result = input_1;
      end
      7'b0000010 : begin
        result = input_2;
      end
      7'b0000011 : begin
        result = input_3;
      end
      7'b0000100 : begin
        result = input_4;
      end
      7'b0000101 : begin
        result = input_5;
      end
      7'b0000110 : begin
        result = input_6;
      end
      7'b0000111 : begin
        result = input_7;
      end
      7'b0001000 : begin
        result = input_8;
      end
      7'b0001001 : begin
        result = input_9;
      end
      7'b0001010 : begin
        result = input_10;
      end
      7'b0001011 : begin
        result = input_11;
      end
      7'b0001100 : begin
        result = input_12;
      end
      7'b0001101 : begin
        result = input_13;
      end
      7'b0001110 : begin
        result = input_14;
      end
      7'b0001111 : begin
        result = input_15;
      end
      7'b0010000 : begin
        result = input_16;
      end
      7'b0010001 : begin
        result = input_17;
      end
      7'b0010010 : begin
        result = input_18;
      end
      7'b0010011 : begin
        result = input_19;
      end
      7'b0010100 : begin
        result = input_20;
      end
      7'b0010101 : begin
        result = input_21;
      end
      7'b0010110 : begin
        result = input_22;
      end
      7'b0010111 : begin
        result = input_23;
      end
      7'b0011000 : begin
        result = input_24;
      end
      7'b0011001 : begin
        result = input_25;
      end
      7'b0011010 : begin
        result = input_26;
      end
      7'b0011011 : begin
        result = input_27;
      end
      7'b0011100 : begin
        result = input_28;
      end
      7'b0011101 : begin
        result = input_29;
      end
      7'b0011110 : begin
        result = input_30;
      end
      7'b0011111 : begin
        result = input_31;
      end
      7'b0100000 : begin
        result = input_32;
      end
      7'b0100001 : begin
        result = input_33;
      end
      7'b0100010 : begin
        result = input_34;
      end
      7'b0100011 : begin
        result = input_35;
      end
      7'b0100100 : begin
        result = input_36;
      end
      7'b0100101 : begin
        result = input_37;
      end
      7'b0100110 : begin
        result = input_38;
      end
      7'b0100111 : begin
        result = input_39;
      end
      7'b0101000 : begin
        result = input_40;
      end
      7'b0101001 : begin
        result = input_41;
      end
      7'b0101010 : begin
        result = input_42;
      end
      7'b0101011 : begin
        result = input_43;
      end
      7'b0101100 : begin
        result = input_44;
      end
      7'b0101101 : begin
        result = input_45;
      end
      7'b0101110 : begin
        result = input_46;
      end
      7'b0101111 : begin
        result = input_47;
      end
      7'b0110000 : begin
        result = input_48;
      end
      7'b0110001 : begin
        result = input_49;
      end
      7'b0110010 : begin
        result = input_50;
      end
      7'b0110011 : begin
        result = input_51;
      end
      7'b0110100 : begin
        result = input_52;
      end
      7'b0110101 : begin
        result = input_53;
      end
      7'b0110110 : begin
        result = input_54;
      end
      7'b0110111 : begin
        result = input_55;
      end
      7'b0111000 : begin
        result = input_56;
      end
      7'b0111001 : begin
        result = input_57;
      end
      7'b0111010 : begin
        result = input_58;
      end
      7'b0111011 : begin
        result = input_59;
      end
      7'b0111100 : begin
        result = input_60;
      end
      7'b0111101 : begin
        result = input_61;
      end
      7'b0111110 : begin
        result = input_62;
      end
      7'b0111111 : begin
        result = input_63;
      end
      7'b1000000 : begin
        result = input_64;
      end
      7'b1000001 : begin
        result = input_65;
      end
      7'b1000010 : begin
        result = input_66;
      end
      7'b1000011 : begin
        result = input_67;
      end
      7'b1000100 : begin
        result = input_68;
      end
      7'b1000101 : begin
        result = input_69;
      end
      7'b1000110 : begin
        result = input_70;
      end
      7'b1000111 : begin
        result = input_71;
      end
      7'b1001000 : begin
        result = input_72;
      end
      7'b1001001 : begin
        result = input_73;
      end
      7'b1001010 : begin
        result = input_74;
      end
      7'b1001011 : begin
        result = input_75;
      end
      7'b1001100 : begin
        result = input_76;
      end
      7'b1001101 : begin
        result = input_77;
      end
      7'b1001110 : begin
        result = input_78;
      end
      7'b1001111 : begin
        result = input_79;
      end
      7'b1010000 : begin
        result = input_80;
      end
      7'b1010001 : begin
        result = input_81;
      end
      7'b1010010 : begin
        result = input_82;
      end
      7'b1010011 : begin
        result = input_83;
      end
      7'b1010100 : begin
        result = input_84;
      end
      7'b1010101 : begin
        result = input_85;
      end
      7'b1010110 : begin
        result = input_86;
      end
      7'b1010111 : begin
        result = input_87;
      end
      7'b1011000 : begin
        result = input_88;
      end
      7'b1011001 : begin
        result = input_89;
      end
      7'b1011010 : begin
        result = input_90;
      end
      7'b1011011 : begin
        result = input_91;
      end
      7'b1011100 : begin
        result = input_92;
      end
      7'b1011101 : begin
        result = input_93;
      end
      7'b1011110 : begin
        result = input_94;
      end
      7'b1011111 : begin
        result = input_95;
      end
      7'b1100000 : begin
        result = input_96;
      end
      7'b1100001 : begin
        result = input_97;
      end
      7'b1100010 : begin
        result = input_98;
      end
      7'b1100011 : begin
        result = input_99;
      end
      7'b1100100 : begin
        result = input_100;
      end
      7'b1100101 : begin
        result = input_101;
      end
      7'b1100110 : begin
        result = input_102;
      end
      7'b1100111 : begin
        result = input_103;
      end
      7'b1101000 : begin
        result = input_104;
      end
      7'b1101001 : begin
        result = input_105;
      end
      7'b1101010 : begin
        result = input_106;
      end
      7'b1101011 : begin
        result = input_107;
      end
      7'b1101100 : begin
        result = input_108;
      end
      7'b1101101 : begin
        result = input_109;
      end
      7'b1101110 : begin
        result = input_110;
      end
      7'b1101111 : begin
        result = input_111;
      end
      7'b1110000 : begin
        result = input_112;
      end
      7'b1110001 : begin
        result = input_113;
      end
      7'b1110010 : begin
        result = input_114;
      end
      7'b1110011 : begin
        result = input_115;
      end
      7'b1110100 : begin
        result = input_116;
      end
      7'b1110101 : begin
        result = input_117;
      end
      7'b1110110 : begin
        result = input_118;
      end
      7'b1110111 : begin
        result = input_119;
      end
      7'b1111000 : begin
        result = input_120;
      end
      7'b1111001 : begin
        result = input_121;
      end
      7'b1111010 : begin
        result = input_122;
      end
      7'b1111011 : begin
        result = input_123;
      end
      7'b1111100 : begin
        result = input_124;
      end
      7'b1111101 : begin
        result = input_125;
      end
      default : begin
        result = input_126;
      end
    endcase
    MUX_v_10_127_2 = result;
  end
  endfunction


  function automatic [12:0] MUX_v_13_2_2;
    input [12:0] input_0;
    input [12:0] input_1;
    input [0:0] sel;
    reg [12:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_13_2_2 = result;
  end
  endfunction


  function automatic [18:0] MUX_v_19_2_2;
    input [18:0] input_0;
    input [18:0] input_1;
    input [0:0] sel;
    reg [18:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_19_2_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input [0:0] sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_127_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [2:0] input_4;
    input [2:0] input_5;
    input [2:0] input_6;
    input [2:0] input_7;
    input [2:0] input_8;
    input [2:0] input_9;
    input [2:0] input_10;
    input [2:0] input_11;
    input [2:0] input_12;
    input [2:0] input_13;
    input [2:0] input_14;
    input [2:0] input_15;
    input [2:0] input_16;
    input [2:0] input_17;
    input [2:0] input_18;
    input [2:0] input_19;
    input [2:0] input_20;
    input [2:0] input_21;
    input [2:0] input_22;
    input [2:0] input_23;
    input [2:0] input_24;
    input [2:0] input_25;
    input [2:0] input_26;
    input [2:0] input_27;
    input [2:0] input_28;
    input [2:0] input_29;
    input [2:0] input_30;
    input [2:0] input_31;
    input [2:0] input_32;
    input [2:0] input_33;
    input [2:0] input_34;
    input [2:0] input_35;
    input [2:0] input_36;
    input [2:0] input_37;
    input [2:0] input_38;
    input [2:0] input_39;
    input [2:0] input_40;
    input [2:0] input_41;
    input [2:0] input_42;
    input [2:0] input_43;
    input [2:0] input_44;
    input [2:0] input_45;
    input [2:0] input_46;
    input [2:0] input_47;
    input [2:0] input_48;
    input [2:0] input_49;
    input [2:0] input_50;
    input [2:0] input_51;
    input [2:0] input_52;
    input [2:0] input_53;
    input [2:0] input_54;
    input [2:0] input_55;
    input [2:0] input_56;
    input [2:0] input_57;
    input [2:0] input_58;
    input [2:0] input_59;
    input [2:0] input_60;
    input [2:0] input_61;
    input [2:0] input_62;
    input [2:0] input_63;
    input [2:0] input_64;
    input [2:0] input_65;
    input [2:0] input_66;
    input [2:0] input_67;
    input [2:0] input_68;
    input [2:0] input_69;
    input [2:0] input_70;
    input [2:0] input_71;
    input [2:0] input_72;
    input [2:0] input_73;
    input [2:0] input_74;
    input [2:0] input_75;
    input [2:0] input_76;
    input [2:0] input_77;
    input [2:0] input_78;
    input [2:0] input_79;
    input [2:0] input_80;
    input [2:0] input_81;
    input [2:0] input_82;
    input [2:0] input_83;
    input [2:0] input_84;
    input [2:0] input_85;
    input [2:0] input_86;
    input [2:0] input_87;
    input [2:0] input_88;
    input [2:0] input_89;
    input [2:0] input_90;
    input [2:0] input_91;
    input [2:0] input_92;
    input [2:0] input_93;
    input [2:0] input_94;
    input [2:0] input_95;
    input [2:0] input_96;
    input [2:0] input_97;
    input [2:0] input_98;
    input [2:0] input_99;
    input [2:0] input_100;
    input [2:0] input_101;
    input [2:0] input_102;
    input [2:0] input_103;
    input [2:0] input_104;
    input [2:0] input_105;
    input [2:0] input_106;
    input [2:0] input_107;
    input [2:0] input_108;
    input [2:0] input_109;
    input [2:0] input_110;
    input [2:0] input_111;
    input [2:0] input_112;
    input [2:0] input_113;
    input [2:0] input_114;
    input [2:0] input_115;
    input [2:0] input_116;
    input [2:0] input_117;
    input [2:0] input_118;
    input [2:0] input_119;
    input [2:0] input_120;
    input [2:0] input_121;
    input [2:0] input_122;
    input [2:0] input_123;
    input [2:0] input_124;
    input [2:0] input_125;
    input [2:0] input_126;
    input [6:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      7'b0000000 : begin
        result = input_0;
      end
      7'b0000001 : begin
        result = input_1;
      end
      7'b0000010 : begin
        result = input_2;
      end
      7'b0000011 : begin
        result = input_3;
      end
      7'b0000100 : begin
        result = input_4;
      end
      7'b0000101 : begin
        result = input_5;
      end
      7'b0000110 : begin
        result = input_6;
      end
      7'b0000111 : begin
        result = input_7;
      end
      7'b0001000 : begin
        result = input_8;
      end
      7'b0001001 : begin
        result = input_9;
      end
      7'b0001010 : begin
        result = input_10;
      end
      7'b0001011 : begin
        result = input_11;
      end
      7'b0001100 : begin
        result = input_12;
      end
      7'b0001101 : begin
        result = input_13;
      end
      7'b0001110 : begin
        result = input_14;
      end
      7'b0001111 : begin
        result = input_15;
      end
      7'b0010000 : begin
        result = input_16;
      end
      7'b0010001 : begin
        result = input_17;
      end
      7'b0010010 : begin
        result = input_18;
      end
      7'b0010011 : begin
        result = input_19;
      end
      7'b0010100 : begin
        result = input_20;
      end
      7'b0010101 : begin
        result = input_21;
      end
      7'b0010110 : begin
        result = input_22;
      end
      7'b0010111 : begin
        result = input_23;
      end
      7'b0011000 : begin
        result = input_24;
      end
      7'b0011001 : begin
        result = input_25;
      end
      7'b0011010 : begin
        result = input_26;
      end
      7'b0011011 : begin
        result = input_27;
      end
      7'b0011100 : begin
        result = input_28;
      end
      7'b0011101 : begin
        result = input_29;
      end
      7'b0011110 : begin
        result = input_30;
      end
      7'b0011111 : begin
        result = input_31;
      end
      7'b0100000 : begin
        result = input_32;
      end
      7'b0100001 : begin
        result = input_33;
      end
      7'b0100010 : begin
        result = input_34;
      end
      7'b0100011 : begin
        result = input_35;
      end
      7'b0100100 : begin
        result = input_36;
      end
      7'b0100101 : begin
        result = input_37;
      end
      7'b0100110 : begin
        result = input_38;
      end
      7'b0100111 : begin
        result = input_39;
      end
      7'b0101000 : begin
        result = input_40;
      end
      7'b0101001 : begin
        result = input_41;
      end
      7'b0101010 : begin
        result = input_42;
      end
      7'b0101011 : begin
        result = input_43;
      end
      7'b0101100 : begin
        result = input_44;
      end
      7'b0101101 : begin
        result = input_45;
      end
      7'b0101110 : begin
        result = input_46;
      end
      7'b0101111 : begin
        result = input_47;
      end
      7'b0110000 : begin
        result = input_48;
      end
      7'b0110001 : begin
        result = input_49;
      end
      7'b0110010 : begin
        result = input_50;
      end
      7'b0110011 : begin
        result = input_51;
      end
      7'b0110100 : begin
        result = input_52;
      end
      7'b0110101 : begin
        result = input_53;
      end
      7'b0110110 : begin
        result = input_54;
      end
      7'b0110111 : begin
        result = input_55;
      end
      7'b0111000 : begin
        result = input_56;
      end
      7'b0111001 : begin
        result = input_57;
      end
      7'b0111010 : begin
        result = input_58;
      end
      7'b0111011 : begin
        result = input_59;
      end
      7'b0111100 : begin
        result = input_60;
      end
      7'b0111101 : begin
        result = input_61;
      end
      7'b0111110 : begin
        result = input_62;
      end
      7'b0111111 : begin
        result = input_63;
      end
      7'b1000000 : begin
        result = input_64;
      end
      7'b1000001 : begin
        result = input_65;
      end
      7'b1000010 : begin
        result = input_66;
      end
      7'b1000011 : begin
        result = input_67;
      end
      7'b1000100 : begin
        result = input_68;
      end
      7'b1000101 : begin
        result = input_69;
      end
      7'b1000110 : begin
        result = input_70;
      end
      7'b1000111 : begin
        result = input_71;
      end
      7'b1001000 : begin
        result = input_72;
      end
      7'b1001001 : begin
        result = input_73;
      end
      7'b1001010 : begin
        result = input_74;
      end
      7'b1001011 : begin
        result = input_75;
      end
      7'b1001100 : begin
        result = input_76;
      end
      7'b1001101 : begin
        result = input_77;
      end
      7'b1001110 : begin
        result = input_78;
      end
      7'b1001111 : begin
        result = input_79;
      end
      7'b1010000 : begin
        result = input_80;
      end
      7'b1010001 : begin
        result = input_81;
      end
      7'b1010010 : begin
        result = input_82;
      end
      7'b1010011 : begin
        result = input_83;
      end
      7'b1010100 : begin
        result = input_84;
      end
      7'b1010101 : begin
        result = input_85;
      end
      7'b1010110 : begin
        result = input_86;
      end
      7'b1010111 : begin
        result = input_87;
      end
      7'b1011000 : begin
        result = input_88;
      end
      7'b1011001 : begin
        result = input_89;
      end
      7'b1011010 : begin
        result = input_90;
      end
      7'b1011011 : begin
        result = input_91;
      end
      7'b1011100 : begin
        result = input_92;
      end
      7'b1011101 : begin
        result = input_93;
      end
      7'b1011110 : begin
        result = input_94;
      end
      7'b1011111 : begin
        result = input_95;
      end
      7'b1100000 : begin
        result = input_96;
      end
      7'b1100001 : begin
        result = input_97;
      end
      7'b1100010 : begin
        result = input_98;
      end
      7'b1100011 : begin
        result = input_99;
      end
      7'b1100100 : begin
        result = input_100;
      end
      7'b1100101 : begin
        result = input_101;
      end
      7'b1100110 : begin
        result = input_102;
      end
      7'b1100111 : begin
        result = input_103;
      end
      7'b1101000 : begin
        result = input_104;
      end
      7'b1101001 : begin
        result = input_105;
      end
      7'b1101010 : begin
        result = input_106;
      end
      7'b1101011 : begin
        result = input_107;
      end
      7'b1101100 : begin
        result = input_108;
      end
      7'b1101101 : begin
        result = input_109;
      end
      7'b1101110 : begin
        result = input_110;
      end
      7'b1101111 : begin
        result = input_111;
      end
      7'b1110000 : begin
        result = input_112;
      end
      7'b1110001 : begin
        result = input_113;
      end
      7'b1110010 : begin
        result = input_114;
      end
      7'b1110011 : begin
        result = input_115;
      end
      7'b1110100 : begin
        result = input_116;
      end
      7'b1110101 : begin
        result = input_117;
      end
      7'b1110110 : begin
        result = input_118;
      end
      7'b1110111 : begin
        result = input_119;
      end
      7'b1111000 : begin
        result = input_120;
      end
      7'b1111001 : begin
        result = input_121;
      end
      7'b1111010 : begin
        result = input_122;
      end
      7'b1111011 : begin
        result = input_123;
      end
      7'b1111100 : begin
        result = input_124;
      end
      7'b1111101 : begin
        result = input_125;
      end
      default : begin
        result = input_126;
      end
    endcase
    MUX_v_3_127_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function automatic [18:0] signext_19_14;
    input [13:0] vector;
  begin
    signext_19_14= {{5{vector[13]}}, vector};
  end
  endfunction


  function automatic [6:0] conv_s2u_2_7 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_7 = {{5{vector[1]}}, vector};
  end
  endfunction


  function automatic [12:0] conv_s2u_13_13 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_13 = vector;
  end
  endfunction


  function automatic [19:0] conv_s2u_13_20 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_20 = {{7{vector[12]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_filter
// ------------------------------------------------------------------


module fir_filter (
  clk, rst, i_sample_rsc_dat, i_sample_rsc_triosy_lz, b_rsc_dat, b_rsc_triosy_lz,
      y_rsc_dat, y_rsc_triosy_lz
);
  input clk;
  input rst;
  input [2:0] i_sample_rsc_dat;
  output i_sample_rsc_triosy_lz;
  input [1269:0] b_rsc_dat;
  output b_rsc_triosy_lz;
  output [8:0] y_rsc_dat;
  output y_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  fir_filter_core fir_filter_core_inst (
      .clk(clk),
      .rst(rst),
      .i_sample_rsc_dat(i_sample_rsc_dat),
      .i_sample_rsc_triosy_lz(i_sample_rsc_triosy_lz),
      .b_rsc_dat(b_rsc_dat),
      .b_rsc_triosy_lz(b_rsc_triosy_lz),
      .y_rsc_dat(y_rsc_dat),
      .y_rsc_triosy_lz(y_rsc_triosy_lz)
    );
endmodule



